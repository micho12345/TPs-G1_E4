module SineWaveLUT (
    input wire [14:0] address,
    output reg [15:0] data
);
    always @(*) begin
        case (address)
            15'b000000000000000 : data = 16'b1000000000000000;
            15'b000000000000001 : data = 16'b1000000000010100;
            15'b000000000000010 : data = 16'b1000000000101001;
            15'b000000000000011 : data = 16'b1000000000111101;
            15'b000000000000100 : data = 16'b1000000001010010;
            15'b000000000000101 : data = 16'b1000000001100110;
            15'b000000000000110 : data = 16'b1000000001111011;
            15'b000000000000111 : data = 16'b1000000010010000;
            15'b000000000001000 : data = 16'b1000000010100100;
            15'b000000000001001 : data = 16'b1000000010111001;
            15'b000000000001010 : data = 16'b1000000011001101;
            15'b000000000001011 : data = 16'b1000000011100010;
            15'b000000000001100 : data = 16'b1000000011110111;
            15'b000000000001101 : data = 16'b1000000100001011;
            15'b000000000001110 : data = 16'b1000000100100000;
            15'b000000000001111 : data = 16'b1000000100110100;
            15'b000000000010000 : data = 16'b1000000101001001;
            15'b000000000010001 : data = 16'b1000000101011101;
            15'b000000000010010 : data = 16'b1000000101110010;
            15'b000000000010011 : data = 16'b1000000110000111;
            15'b000000000010100 : data = 16'b1000000110011011;
            15'b000000000010101 : data = 16'b1000000110110000;
            15'b000000000010110 : data = 16'b1000000111000100;
            15'b000000000010111 : data = 16'b1000000111011001;
            15'b000000000011000 : data = 16'b1000000111101110;
            15'b000000000011001 : data = 16'b1000001000000010;
            15'b000000000011010 : data = 16'b1000001000010111;
            15'b000000000011011 : data = 16'b1000001000101011;
            15'b000000000011100 : data = 16'b1000001001000000;
            15'b000000000011101 : data = 16'b1000001001010101;
            15'b000000000011110 : data = 16'b1000001001101001;
            15'b000000000011111 : data = 16'b1000001001111110;
            15'b000000000100000 : data = 16'b1000001010010010;
            15'b000000000100001 : data = 16'b1000001010100111;
            15'b000000000100010 : data = 16'b1000001010111011;
            15'b000000000100011 : data = 16'b1000001011010000;
            15'b000000000100100 : data = 16'b1000001011100101;
            15'b000000000100101 : data = 16'b1000001011111001;
            15'b000000000100110 : data = 16'b1000001100001110;
            15'b000000000100111 : data = 16'b1000001100100010;
            15'b000000000101000 : data = 16'b1000001100110111;
            15'b000000000101001 : data = 16'b1000001101001100;
            15'b000000000101010 : data = 16'b1000001101100000;
            15'b000000000101011 : data = 16'b1000001101110101;
            15'b000000000101100 : data = 16'b1000001110001001;
            15'b000000000101101 : data = 16'b1000001110011110;
            15'b000000000101110 : data = 16'b1000001110110010;
            15'b000000000101111 : data = 16'b1000001111000111;
            15'b000000000110000 : data = 16'b1000001111011100;
            15'b000000000110001 : data = 16'b1000001111110000;
            15'b000000000110010 : data = 16'b1000010000000101;
            15'b000000000110011 : data = 16'b1000010000011001;
            15'b000000000110100 : data = 16'b1000010000101110;
            15'b000000000110101 : data = 16'b1000010001000010;
            15'b000000000110110 : data = 16'b1000010001010111;
            15'b000000000110111 : data = 16'b1000010001101100;
            15'b000000000111000 : data = 16'b1000010010000000;
            15'b000000000111001 : data = 16'b1000010010010101;
            15'b000000000111010 : data = 16'b1000010010101001;
            15'b000000000111011 : data = 16'b1000010010111110;
            15'b000000000111100 : data = 16'b1000010011010010;
            15'b000000000111101 : data = 16'b1000010011100111;
            15'b000000000111110 : data = 16'b1000010011111100;
            15'b000000000111111 : data = 16'b1000010100010000;
            15'b000000001000000 : data = 16'b1000010100100101;
            15'b000000001000001 : data = 16'b1000010100111001;
            15'b000000001000010 : data = 16'b1000010101001110;
            15'b000000001000011 : data = 16'b1000010101100010;
            15'b000000001000100 : data = 16'b1000010101110111;
            15'b000000001000101 : data = 16'b1000010110001100;
            15'b000000001000110 : data = 16'b1000010110100000;
            15'b000000001000111 : data = 16'b1000010110110101;
            15'b000000001001000 : data = 16'b1000010111001001;
            15'b000000001001001 : data = 16'b1000010111011110;
            15'b000000001001010 : data = 16'b1000010111110010;
            15'b000000001001011 : data = 16'b1000011000000111;
            15'b000000001001100 : data = 16'b1000011000011100;
            15'b000000001001101 : data = 16'b1000011000110000;
            15'b000000001001110 : data = 16'b1000011001000101;
            15'b000000001001111 : data = 16'b1000011001011001;
            15'b000000001010000 : data = 16'b1000011001101110;
            15'b000000001010001 : data = 16'b1000011010000010;
            15'b000000001010010 : data = 16'b1000011010010111;
            15'b000000001010011 : data = 16'b1000011010101100;
            15'b000000001010100 : data = 16'b1000011011000000;
            15'b000000001010101 : data = 16'b1000011011010101;
            15'b000000001010110 : data = 16'b1000011011101001;
            15'b000000001010111 : data = 16'b1000011011111110;
            15'b000000001011000 : data = 16'b1000011100010010;
            15'b000000001011001 : data = 16'b1000011100100111;
            15'b000000001011010 : data = 16'b1000011100111011;
            15'b000000001011011 : data = 16'b1000011101010000;
            15'b000000001011100 : data = 16'b1000011101100101;
            15'b000000001011101 : data = 16'b1000011101111001;
            15'b000000001011110 : data = 16'b1000011110001110;
            15'b000000001011111 : data = 16'b1000011110100010;
            15'b000000001100000 : data = 16'b1000011110110111;
            15'b000000001100001 : data = 16'b1000011111001011;
            15'b000000001100010 : data = 16'b1000011111100000;
            15'b000000001100011 : data = 16'b1000011111110100;
            15'b000000001100100 : data = 16'b1000100000001001;
            15'b000000001100101 : data = 16'b1000100000011110;
            15'b000000001100110 : data = 16'b1000100000110010;
            15'b000000001100111 : data = 16'b1000100001000111;
            15'b000000001101000 : data = 16'b1000100001011011;
            15'b000000001101001 : data = 16'b1000100001110000;
            15'b000000001101010 : data = 16'b1000100010000100;
            15'b000000001101011 : data = 16'b1000100010011001;
            15'b000000001101100 : data = 16'b1000100010101101;
            15'b000000001101101 : data = 16'b1000100011000010;
            15'b000000001101110 : data = 16'b1000100011010110;
            15'b000000001101111 : data = 16'b1000100011101011;
            15'b000000001110000 : data = 16'b1000100011111111;
            15'b000000001110001 : data = 16'b1000100100010100;
            15'b000000001110010 : data = 16'b1000100100101001;
            15'b000000001110011 : data = 16'b1000100100111101;
            15'b000000001110100 : data = 16'b1000100101010010;
            15'b000000001110101 : data = 16'b1000100101100110;
            15'b000000001110110 : data = 16'b1000100101111011;
            15'b000000001110111 : data = 16'b1000100110001111;
            15'b000000001111000 : data = 16'b1000100110100100;
            15'b000000001111001 : data = 16'b1000100110111000;
            15'b000000001111010 : data = 16'b1000100111001101;
            15'b000000001111011 : data = 16'b1000100111100001;
            15'b000000001111100 : data = 16'b1000100111110110;
            15'b000000001111101 : data = 16'b1000101000001010;
            15'b000000001111110 : data = 16'b1000101000011111;
            15'b000000001111111 : data = 16'b1000101000110011;
            15'b000000010000000 : data = 16'b1000101001001000;
            15'b000000010000001 : data = 16'b1000101001011100;
            15'b000000010000010 : data = 16'b1000101001110001;
            15'b000000010000011 : data = 16'b1000101010000101;
            15'b000000010000100 : data = 16'b1000101010011010;
            15'b000000010000101 : data = 16'b1000101010101111;
            15'b000000010000110 : data = 16'b1000101011000011;
            15'b000000010000111 : data = 16'b1000101011011000;
            15'b000000010001000 : data = 16'b1000101011101100;
            15'b000000010001001 : data = 16'b1000101100000001;
            15'b000000010001010 : data = 16'b1000101100010101;
            15'b000000010001011 : data = 16'b1000101100101010;
            15'b000000010001100 : data = 16'b1000101100111110;
            15'b000000010001101 : data = 16'b1000101101010011;
            15'b000000010001110 : data = 16'b1000101101100111;
            15'b000000010001111 : data = 16'b1000101101111100;
            15'b000000010010000 : data = 16'b1000101110010000;
            15'b000000010010001 : data = 16'b1000101110100101;
            15'b000000010010010 : data = 16'b1000101110111001;
            15'b000000010010011 : data = 16'b1000101111001110;
            15'b000000010010100 : data = 16'b1000101111100010;
            15'b000000010010101 : data = 16'b1000101111110111;
            15'b000000010010110 : data = 16'b1000110000001011;
            15'b000000010010111 : data = 16'b1000110000100000;
            15'b000000010011000 : data = 16'b1000110000110100;
            15'b000000010011001 : data = 16'b1000110001001001;
            15'b000000010011010 : data = 16'b1000110001011101;
            15'b000000010011011 : data = 16'b1000110001110010;
            15'b000000010011100 : data = 16'b1000110010000110;
            15'b000000010011101 : data = 16'b1000110010011011;
            15'b000000010011110 : data = 16'b1000110010101111;
            15'b000000010011111 : data = 16'b1000110011000100;
            15'b000000010100000 : data = 16'b1000110011011000;
            15'b000000010100001 : data = 16'b1000110011101101;
            15'b000000010100010 : data = 16'b1000110100000001;
            15'b000000010100011 : data = 16'b1000110100010101;
            15'b000000010100100 : data = 16'b1000110100101010;
            15'b000000010100101 : data = 16'b1000110100111110;
            15'b000000010100110 : data = 16'b1000110101010011;
            15'b000000010100111 : data = 16'b1000110101100111;
            15'b000000010101000 : data = 16'b1000110101111100;
            15'b000000010101001 : data = 16'b1000110110010000;
            15'b000000010101010 : data = 16'b1000110110100101;
            15'b000000010101011 : data = 16'b1000110110111001;
            15'b000000010101100 : data = 16'b1000110111001110;
            15'b000000010101101 : data = 16'b1000110111100010;
            15'b000000010101110 : data = 16'b1000110111110111;
            15'b000000010101111 : data = 16'b1000111000001011;
            15'b000000010110000 : data = 16'b1000111000100000;
            15'b000000010110001 : data = 16'b1000111000110100;
            15'b000000010110010 : data = 16'b1000111001001001;
            15'b000000010110011 : data = 16'b1000111001011101;
            15'b000000010110100 : data = 16'b1000111001110001;
            15'b000000010110101 : data = 16'b1000111010000110;
            15'b000000010110110 : data = 16'b1000111010011010;
            15'b000000010110111 : data = 16'b1000111010101111;
            15'b000000010111000 : data = 16'b1000111011000011;
            15'b000000010111001 : data = 16'b1000111011011000;
            15'b000000010111010 : data = 16'b1000111011101100;
            15'b000000010111011 : data = 16'b1000111100000001;
            15'b000000010111100 : data = 16'b1000111100010101;
            15'b000000010111101 : data = 16'b1000111100101010;
            15'b000000010111110 : data = 16'b1000111100111110;
            15'b000000010111111 : data = 16'b1000111101010010;
            15'b000000011000000 : data = 16'b1000111101100111;
            15'b000000011000001 : data = 16'b1000111101111011;
            15'b000000011000010 : data = 16'b1000111110010000;
            15'b000000011000011 : data = 16'b1000111110100100;
            15'b000000011000100 : data = 16'b1000111110111001;
            15'b000000011000101 : data = 16'b1000111111001101;
            15'b000000011000110 : data = 16'b1000111111100001;
            15'b000000011000111 : data = 16'b1000111111110110;
            15'b000000011001000 : data = 16'b1001000000001010;
            15'b000000011001001 : data = 16'b1001000000011111;
            15'b000000011001010 : data = 16'b1001000000110011;
            15'b000000011001011 : data = 16'b1001000001001000;
            15'b000000011001100 : data = 16'b1001000001011100;
            15'b000000011001101 : data = 16'b1001000001110000;
            15'b000000011001110 : data = 16'b1001000010000101;
            15'b000000011001111 : data = 16'b1001000010011001;
            15'b000000011010000 : data = 16'b1001000010101110;
            15'b000000011010001 : data = 16'b1001000011000010;
            15'b000000011010010 : data = 16'b1001000011010110;
            15'b000000011010011 : data = 16'b1001000011101011;
            15'b000000011010100 : data = 16'b1001000011111111;
            15'b000000011010101 : data = 16'b1001000100010100;
            15'b000000011010110 : data = 16'b1001000100101000;
            15'b000000011010111 : data = 16'b1001000100111100;
            15'b000000011011000 : data = 16'b1001000101010001;
            15'b000000011011001 : data = 16'b1001000101100101;
            15'b000000011011010 : data = 16'b1001000101111010;
            15'b000000011011011 : data = 16'b1001000110001110;
            15'b000000011011100 : data = 16'b1001000110100010;
            15'b000000011011101 : data = 16'b1001000110110111;
            15'b000000011011110 : data = 16'b1001000111001011;
            15'b000000011011111 : data = 16'b1001000111100000;
            15'b000000011100000 : data = 16'b1001000111110100;
            15'b000000011100001 : data = 16'b1001001000001000;
            15'b000000011100010 : data = 16'b1001001000011101;
            15'b000000011100011 : data = 16'b1001001000110001;
            15'b000000011100100 : data = 16'b1001001001000110;
            15'b000000011100101 : data = 16'b1001001001011010;
            15'b000000011100110 : data = 16'b1001001001101110;
            15'b000000011100111 : data = 16'b1001001010000011;
            15'b000000011101000 : data = 16'b1001001010010111;
            15'b000000011101001 : data = 16'b1001001010101011;
            15'b000000011101010 : data = 16'b1001001011000000;
            15'b000000011101011 : data = 16'b1001001011010100;
            15'b000000011101100 : data = 16'b1001001011101001;
            15'b000000011101101 : data = 16'b1001001011111101;
            15'b000000011101110 : data = 16'b1001001100010001;
            15'b000000011101111 : data = 16'b1001001100100110;
            15'b000000011110000 : data = 16'b1001001100111010;
            15'b000000011110001 : data = 16'b1001001101001110;
            15'b000000011110010 : data = 16'b1001001101100011;
            15'b000000011110011 : data = 16'b1001001101110111;
            15'b000000011110100 : data = 16'b1001001110001011;
            15'b000000011110101 : data = 16'b1001001110100000;
            15'b000000011110110 : data = 16'b1001001110110100;
            15'b000000011110111 : data = 16'b1001001111001000;
            15'b000000011111000 : data = 16'b1001001111011101;
            15'b000000011111001 : data = 16'b1001001111110001;
            15'b000000011111010 : data = 16'b1001010000000101;
            15'b000000011111011 : data = 16'b1001010000011010;
            15'b000000011111100 : data = 16'b1001010000101110;
            15'b000000011111101 : data = 16'b1001010001000010;
            15'b000000011111110 : data = 16'b1001010001010111;
            15'b000000011111111 : data = 16'b1001010001101011;
            15'b000000100000000 : data = 16'b1001010001111111;
            15'b000000100000001 : data = 16'b1001010010010100;
            15'b000000100000010 : data = 16'b1001010010101000;
            15'b000000100000011 : data = 16'b1001010010111100;
            15'b000000100000100 : data = 16'b1001010011010001;
            15'b000000100000101 : data = 16'b1001010011100101;
            15'b000000100000110 : data = 16'b1001010011111001;
            15'b000000100000111 : data = 16'b1001010100001110;
            15'b000000100001000 : data = 16'b1001010100100010;
            15'b000000100001001 : data = 16'b1001010100110110;
            15'b000000100001010 : data = 16'b1001010101001010;
            15'b000000100001011 : data = 16'b1001010101011111;
            15'b000000100001100 : data = 16'b1001010101110011;
            15'b000000100001101 : data = 16'b1001010110000111;
            15'b000000100001110 : data = 16'b1001010110011100;
            15'b000000100001111 : data = 16'b1001010110110000;
            15'b000000100010000 : data = 16'b1001010111000100;
            15'b000000100010001 : data = 16'b1001010111011001;
            15'b000000100010010 : data = 16'b1001010111101101;
            15'b000000100010011 : data = 16'b1001011000000001;
            15'b000000100010100 : data = 16'b1001011000010101;
            15'b000000100010101 : data = 16'b1001011000101010;
            15'b000000100010110 : data = 16'b1001011000111110;
            15'b000000100010111 : data = 16'b1001011001010010;
            15'b000000100011000 : data = 16'b1001011001100110;
            15'b000000100011001 : data = 16'b1001011001111011;
            15'b000000100011010 : data = 16'b1001011010001111;
            15'b000000100011011 : data = 16'b1001011010100011;
            15'b000000100011100 : data = 16'b1001011010111000;
            15'b000000100011101 : data = 16'b1001011011001100;
            15'b000000100011110 : data = 16'b1001011011100000;
            15'b000000100011111 : data = 16'b1001011011110100;
            15'b000000100100000 : data = 16'b1001011100001001;
            15'b000000100100001 : data = 16'b1001011100011101;
            15'b000000100100010 : data = 16'b1001011100110001;
            15'b000000100100011 : data = 16'b1001011101000101;
            15'b000000100100100 : data = 16'b1001011101011010;
            15'b000000100100101 : data = 16'b1001011101101110;
            15'b000000100100110 : data = 16'b1001011110000010;
            15'b000000100100111 : data = 16'b1001011110010110;
            15'b000000100101000 : data = 16'b1001011110101011;
            15'b000000100101001 : data = 16'b1001011110111111;
            15'b000000100101010 : data = 16'b1001011111010011;
            15'b000000100101011 : data = 16'b1001011111100111;
            15'b000000100101100 : data = 16'b1001011111111011;
            15'b000000100101101 : data = 16'b1001100000010000;
            15'b000000100101110 : data = 16'b1001100000100100;
            15'b000000100101111 : data = 16'b1001100000111000;
            15'b000000100110000 : data = 16'b1001100001001100;
            15'b000000100110001 : data = 16'b1001100001100001;
            15'b000000100110010 : data = 16'b1001100001110101;
            15'b000000100110011 : data = 16'b1001100010001001;
            15'b000000100110100 : data = 16'b1001100010011101;
            15'b000000100110101 : data = 16'b1001100010110001;
            15'b000000100110110 : data = 16'b1001100011000110;
            15'b000000100110111 : data = 16'b1001100011011010;
            15'b000000100111000 : data = 16'b1001100011101110;
            15'b000000100111001 : data = 16'b1001100100000010;
            15'b000000100111010 : data = 16'b1001100100010110;
            15'b000000100111011 : data = 16'b1001100100101010;
            15'b000000100111100 : data = 16'b1001100100111111;
            15'b000000100111101 : data = 16'b1001100101010011;
            15'b000000100111110 : data = 16'b1001100101100111;
            15'b000000100111111 : data = 16'b1001100101111011;
            15'b000000101000000 : data = 16'b1001100110001111;
            15'b000000101000001 : data = 16'b1001100110100100;
            15'b000000101000010 : data = 16'b1001100110111000;
            15'b000000101000011 : data = 16'b1001100111001100;
            15'b000000101000100 : data = 16'b1001100111100000;
            15'b000000101000101 : data = 16'b1001100111110100;
            15'b000000101000110 : data = 16'b1001101000001000;
            15'b000000101000111 : data = 16'b1001101000011101;
            15'b000000101001000 : data = 16'b1001101000110001;
            15'b000000101001001 : data = 16'b1001101001000101;
            15'b000000101001010 : data = 16'b1001101001011001;
            15'b000000101001011 : data = 16'b1001101001101101;
            15'b000000101001100 : data = 16'b1001101010000001;
            15'b000000101001101 : data = 16'b1001101010010101;
            15'b000000101001110 : data = 16'b1001101010101010;
            15'b000000101001111 : data = 16'b1001101010111110;
            15'b000000101010000 : data = 16'b1001101011010010;
            15'b000000101010001 : data = 16'b1001101011100110;
            15'b000000101010010 : data = 16'b1001101011111010;
            15'b000000101010011 : data = 16'b1001101100001110;
            15'b000000101010100 : data = 16'b1001101100100010;
            15'b000000101010101 : data = 16'b1001101100110110;
            15'b000000101010110 : data = 16'b1001101101001011;
            15'b000000101010111 : data = 16'b1001101101011111;
            15'b000000101011000 : data = 16'b1001101101110011;
            15'b000000101011001 : data = 16'b1001101110000111;
            15'b000000101011010 : data = 16'b1001101110011011;
            15'b000000101011011 : data = 16'b1001101110101111;
            15'b000000101011100 : data = 16'b1001101111000011;
            15'b000000101011101 : data = 16'b1001101111010111;
            15'b000000101011110 : data = 16'b1001101111101011;
            15'b000000101011111 : data = 16'b1001101111111111;
            15'b000000101100000 : data = 16'b1001110000010100;
            15'b000000101100001 : data = 16'b1001110000101000;
            15'b000000101100010 : data = 16'b1001110000111100;
            15'b000000101100011 : data = 16'b1001110001010000;
            15'b000000101100100 : data = 16'b1001110001100100;
            15'b000000101100101 : data = 16'b1001110001111000;
            15'b000000101100110 : data = 16'b1001110010001100;
            15'b000000101100111 : data = 16'b1001110010100000;
            15'b000000101101000 : data = 16'b1001110010110100;
            15'b000000101101001 : data = 16'b1001110011001000;
            15'b000000101101010 : data = 16'b1001110011011100;
            15'b000000101101011 : data = 16'b1001110011110000;
            15'b000000101101100 : data = 16'b1001110100000100;
            15'b000000101101101 : data = 16'b1001110100011000;
            15'b000000101101110 : data = 16'b1001110100101101;
            15'b000000101101111 : data = 16'b1001110101000001;
            15'b000000101110000 : data = 16'b1001110101010101;
            15'b000000101110001 : data = 16'b1001110101101001;
            15'b000000101110010 : data = 16'b1001110101111101;
            15'b000000101110011 : data = 16'b1001110110010001;
            15'b000000101110100 : data = 16'b1001110110100101;
            15'b000000101110101 : data = 16'b1001110110111001;
            15'b000000101110110 : data = 16'b1001110111001101;
            15'b000000101110111 : data = 16'b1001110111100001;
            15'b000000101111000 : data = 16'b1001110111110101;
            15'b000000101111001 : data = 16'b1001111000001001;
            15'b000000101111010 : data = 16'b1001111000011101;
            15'b000000101111011 : data = 16'b1001111000110001;
            15'b000000101111100 : data = 16'b1001111001000101;
            15'b000000101111101 : data = 16'b1001111001011001;
            15'b000000101111110 : data = 16'b1001111001101101;
            15'b000000101111111 : data = 16'b1001111010000001;
            15'b000000110000000 : data = 16'b1001111010010101;
            15'b000000110000001 : data = 16'b1001111010101001;
            15'b000000110000010 : data = 16'b1001111010111101;
            15'b000000110000011 : data = 16'b1001111011010001;
            15'b000000110000100 : data = 16'b1001111011100101;
            15'b000000110000101 : data = 16'b1001111011111001;
            15'b000000110000110 : data = 16'b1001111100001101;
            15'b000000110000111 : data = 16'b1001111100100001;
            15'b000000110001000 : data = 16'b1001111100110101;
            15'b000000110001001 : data = 16'b1001111101001001;
            15'b000000110001010 : data = 16'b1001111101011101;
            15'b000000110001011 : data = 16'b1001111101110001;
            15'b000000110001100 : data = 16'b1001111110000101;
            15'b000000110001101 : data = 16'b1001111110011000;
            15'b000000110001110 : data = 16'b1001111110101100;
            15'b000000110001111 : data = 16'b1001111111000000;
            15'b000000110010000 : data = 16'b1001111111010100;
            15'b000000110010001 : data = 16'b1001111111101000;
            15'b000000110010010 : data = 16'b1001111111111100;
            15'b000000110010011 : data = 16'b1010000000010000;
            15'b000000110010100 : data = 16'b1010000000100100;
            15'b000000110010101 : data = 16'b1010000000111000;
            15'b000000110010110 : data = 16'b1010000001001100;
            15'b000000110010111 : data = 16'b1010000001100000;
            15'b000000110011000 : data = 16'b1010000001110100;
            15'b000000110011001 : data = 16'b1010000010001000;
            15'b000000110011010 : data = 16'b1010000010011100;
            15'b000000110011011 : data = 16'b1010000010101111;
            15'b000000110011100 : data = 16'b1010000011000011;
            15'b000000110011101 : data = 16'b1010000011010111;
            15'b000000110011110 : data = 16'b1010000011101011;
            15'b000000110011111 : data = 16'b1010000011111111;
            15'b000000110100000 : data = 16'b1010000100010011;
            15'b000000110100001 : data = 16'b1010000100100111;
            15'b000000110100010 : data = 16'b1010000100111011;
            15'b000000110100011 : data = 16'b1010000101001111;
            15'b000000110100100 : data = 16'b1010000101100010;
            15'b000000110100101 : data = 16'b1010000101110110;
            15'b000000110100110 : data = 16'b1010000110001010;
            15'b000000110100111 : data = 16'b1010000110011110;
            15'b000000110101000 : data = 16'b1010000110110010;
            15'b000000110101001 : data = 16'b1010000111000110;
            15'b000000110101010 : data = 16'b1010000111011010;
            15'b000000110101011 : data = 16'b1010000111101110;
            15'b000000110101100 : data = 16'b1010001000000001;
            15'b000000110101101 : data = 16'b1010001000010101;
            15'b000000110101110 : data = 16'b1010001000101001;
            15'b000000110101111 : data = 16'b1010001000111101;
            15'b000000110110000 : data = 16'b1010001001010001;
            15'b000000110110001 : data = 16'b1010001001100101;
            15'b000000110110010 : data = 16'b1010001001111000;
            15'b000000110110011 : data = 16'b1010001010001100;
            15'b000000110110100 : data = 16'b1010001010100000;
            15'b000000110110101 : data = 16'b1010001010110100;
            15'b000000110110110 : data = 16'b1010001011001000;
            15'b000000110110111 : data = 16'b1010001011011100;
            15'b000000110111000 : data = 16'b1010001011101111;
            15'b000000110111001 : data = 16'b1010001100000011;
            15'b000000110111010 : data = 16'b1010001100010111;
            15'b000000110111011 : data = 16'b1010001100101011;
            15'b000000110111100 : data = 16'b1010001100111111;
            15'b000000110111101 : data = 16'b1010001101010010;
            15'b000000110111110 : data = 16'b1010001101100110;
            15'b000000110111111 : data = 16'b1010001101111010;
            15'b000000111000000 : data = 16'b1010001110001110;
            15'b000000111000001 : data = 16'b1010001110100001;
            15'b000000111000010 : data = 16'b1010001110110101;
            15'b000000111000011 : data = 16'b1010001111001001;
            15'b000000111000100 : data = 16'b1010001111011101;
            15'b000000111000101 : data = 16'b1010001111110000;
            15'b000000111000110 : data = 16'b1010010000000100;
            15'b000000111000111 : data = 16'b1010010000011000;
            15'b000000111001000 : data = 16'b1010010000101100;
            15'b000000111001001 : data = 16'b1010010001000000;
            15'b000000111001010 : data = 16'b1010010001010011;
            15'b000000111001011 : data = 16'b1010010001100111;
            15'b000000111001100 : data = 16'b1010010001111011;
            15'b000000111001101 : data = 16'b1010010010001110;
            15'b000000111001110 : data = 16'b1010010010100010;
            15'b000000111001111 : data = 16'b1010010010110110;
            15'b000000111010000 : data = 16'b1010010011001010;
            15'b000000111010001 : data = 16'b1010010011011101;
            15'b000000111010010 : data = 16'b1010010011110001;
            15'b000000111010011 : data = 16'b1010010100000101;
            15'b000000111010100 : data = 16'b1010010100011000;
            15'b000000111010101 : data = 16'b1010010100101100;
            15'b000000111010110 : data = 16'b1010010101000000;
            15'b000000111010111 : data = 16'b1010010101010100;
            15'b000000111011000 : data = 16'b1010010101100111;
            15'b000000111011001 : data = 16'b1010010101111011;
            15'b000000111011010 : data = 16'b1010010110001111;
            15'b000000111011011 : data = 16'b1010010110100010;
            15'b000000111011100 : data = 16'b1010010110110110;
            15'b000000111011101 : data = 16'b1010010111001010;
            15'b000000111011110 : data = 16'b1010010111011101;
            15'b000000111011111 : data = 16'b1010010111110001;
            15'b000000111100000 : data = 16'b1010011000000101;
            15'b000000111100001 : data = 16'b1010011000011000;
            15'b000000111100010 : data = 16'b1010011000101100;
            15'b000000111100011 : data = 16'b1010011001000000;
            15'b000000111100100 : data = 16'b1010011001010011;
            15'b000000111100101 : data = 16'b1010011001100111;
            15'b000000111100110 : data = 16'b1010011001111011;
            15'b000000111100111 : data = 16'b1010011010001110;
            15'b000000111101000 : data = 16'b1010011010100010;
            15'b000000111101001 : data = 16'b1010011010110101;
            15'b000000111101010 : data = 16'b1010011011001001;
            15'b000000111101011 : data = 16'b1010011011011101;
            15'b000000111101100 : data = 16'b1010011011110000;
            15'b000000111101101 : data = 16'b1010011100000100;
            15'b000000111101110 : data = 16'b1010011100011000;
            15'b000000111101111 : data = 16'b1010011100101011;
            15'b000000111110000 : data = 16'b1010011100111111;
            15'b000000111110001 : data = 16'b1010011101010010;
            15'b000000111110010 : data = 16'b1010011101100110;
            15'b000000111110011 : data = 16'b1010011101111001;
            15'b000000111110100 : data = 16'b1010011110001101;
            15'b000000111110101 : data = 16'b1010011110100001;
            15'b000000111110110 : data = 16'b1010011110110100;
            15'b000000111110111 : data = 16'b1010011111001000;
            15'b000000111111000 : data = 16'b1010011111011011;
            15'b000000111111001 : data = 16'b1010011111101111;
            15'b000000111111010 : data = 16'b1010100000000010;
            15'b000000111111011 : data = 16'b1010100000010110;
            15'b000000111111100 : data = 16'b1010100000101010;
            15'b000000111111101 : data = 16'b1010100000111101;
            15'b000000111111110 : data = 16'b1010100001010001;
            15'b000000111111111 : data = 16'b1010100001100100;
            15'b000001000000000 : data = 16'b1010100001111000;
            15'b000001000000001 : data = 16'b1010100010001011;
            15'b000001000000010 : data = 16'b1010100010011111;
            15'b000001000000011 : data = 16'b1010100010110010;
            15'b000001000000100 : data = 16'b1010100011000110;
            15'b000001000000101 : data = 16'b1010100011011001;
            15'b000001000000110 : data = 16'b1010100011101101;
            15'b000001000000111 : data = 16'b1010100100000000;
            15'b000001000001000 : data = 16'b1010100100010100;
            15'b000001000001001 : data = 16'b1010100100100111;
            15'b000001000001010 : data = 16'b1010100100111011;
            15'b000001000001011 : data = 16'b1010100101001110;
            15'b000001000001100 : data = 16'b1010100101100010;
            15'b000001000001101 : data = 16'b1010100101110101;
            15'b000001000001110 : data = 16'b1010100110001001;
            15'b000001000001111 : data = 16'b1010100110011100;
            15'b000001000010000 : data = 16'b1010100110110000;
            15'b000001000010001 : data = 16'b1010100111000011;
            15'b000001000010010 : data = 16'b1010100111010111;
            15'b000001000010011 : data = 16'b1010100111101010;
            15'b000001000010100 : data = 16'b1010100111111110;
            15'b000001000010101 : data = 16'b1010101000010001;
            15'b000001000010110 : data = 16'b1010101000100100;
            15'b000001000010111 : data = 16'b1010101000111000;
            15'b000001000011000 : data = 16'b1010101001001011;
            15'b000001000011001 : data = 16'b1010101001011111;
            15'b000001000011010 : data = 16'b1010101001110010;
            15'b000001000011011 : data = 16'b1010101010000110;
            15'b000001000011100 : data = 16'b1010101010011001;
            15'b000001000011101 : data = 16'b1010101010101100;
            15'b000001000011110 : data = 16'b1010101011000000;
            15'b000001000011111 : data = 16'b1010101011010011;
            15'b000001000100000 : data = 16'b1010101011100111;
            15'b000001000100001 : data = 16'b1010101011111010;
            15'b000001000100010 : data = 16'b1010101100001101;
            15'b000001000100011 : data = 16'b1010101100100001;
            15'b000001000100100 : data = 16'b1010101100110100;
            15'b000001000100101 : data = 16'b1010101101001000;
            15'b000001000100110 : data = 16'b1010101101011011;
            15'b000001000100111 : data = 16'b1010101101101110;
            15'b000001000101000 : data = 16'b1010101110000010;
            15'b000001000101001 : data = 16'b1010101110010101;
            15'b000001000101010 : data = 16'b1010101110101000;
            15'b000001000101011 : data = 16'b1010101110111100;
            15'b000001000101100 : data = 16'b1010101111001111;
            15'b000001000101101 : data = 16'b1010101111100010;
            15'b000001000101110 : data = 16'b1010101111110110;
            15'b000001000101111 : data = 16'b1010110000001001;
            15'b000001000110000 : data = 16'b1010110000011100;
            15'b000001000110001 : data = 16'b1010110000110000;
            15'b000001000110010 : data = 16'b1010110001000011;
            15'b000001000110011 : data = 16'b1010110001010110;
            15'b000001000110100 : data = 16'b1010110001101010;
            15'b000001000110101 : data = 16'b1010110001111101;
            15'b000001000110110 : data = 16'b1010110010010000;
            15'b000001000110111 : data = 16'b1010110010100100;
            15'b000001000111000 : data = 16'b1010110010110111;
            15'b000001000111001 : data = 16'b1010110011001010;
            15'b000001000111010 : data = 16'b1010110011011101;
            15'b000001000111011 : data = 16'b1010110011110001;
            15'b000001000111100 : data = 16'b1010110100000100;
            15'b000001000111101 : data = 16'b1010110100010111;
            15'b000001000111110 : data = 16'b1010110100101011;
            15'b000001000111111 : data = 16'b1010110100111110;
            15'b000001001000000 : data = 16'b1010110101010001;
            15'b000001001000001 : data = 16'b1010110101100100;
            15'b000001001000010 : data = 16'b1010110101111000;
            15'b000001001000011 : data = 16'b1010110110001011;
            15'b000001001000100 : data = 16'b1010110110011110;
            15'b000001001000101 : data = 16'b1010110110110001;
            15'b000001001000110 : data = 16'b1010110111000101;
            15'b000001001000111 : data = 16'b1010110111011000;
            15'b000001001001000 : data = 16'b1010110111101011;
            15'b000001001001001 : data = 16'b1010110111111110;
            15'b000001001001010 : data = 16'b1010111000010001;
            15'b000001001001011 : data = 16'b1010111000100101;
            15'b000001001001100 : data = 16'b1010111000111000;
            15'b000001001001101 : data = 16'b1010111001001011;
            15'b000001001001110 : data = 16'b1010111001011110;
            15'b000001001001111 : data = 16'b1010111001110001;
            15'b000001001010000 : data = 16'b1010111010000101;
            15'b000001001010001 : data = 16'b1010111010011000;
            15'b000001001010010 : data = 16'b1010111010101011;
            15'b000001001010011 : data = 16'b1010111010111110;
            15'b000001001010100 : data = 16'b1010111011010001;
            15'b000001001010101 : data = 16'b1010111011100100;
            15'b000001001010110 : data = 16'b1010111011111000;
            15'b000001001010111 : data = 16'b1010111100001011;
            15'b000001001011000 : data = 16'b1010111100011110;
            15'b000001001011001 : data = 16'b1010111100110001;
            15'b000001001011010 : data = 16'b1010111101000100;
            15'b000001001011011 : data = 16'b1010111101010111;
            15'b000001001011100 : data = 16'b1010111101101010;
            15'b000001001011101 : data = 16'b1010111101111101;
            15'b000001001011110 : data = 16'b1010111110010001;
            15'b000001001011111 : data = 16'b1010111110100100;
            15'b000001001100000 : data = 16'b1010111110110111;
            15'b000001001100001 : data = 16'b1010111111001010;
            15'b000001001100010 : data = 16'b1010111111011101;
            15'b000001001100011 : data = 16'b1010111111110000;
            15'b000001001100100 : data = 16'b1011000000000011;
            15'b000001001100101 : data = 16'b1011000000010110;
            15'b000001001100110 : data = 16'b1011000000101001;
            15'b000001001100111 : data = 16'b1011000000111100;
            15'b000001001101000 : data = 16'b1011000001010000;
            15'b000001001101001 : data = 16'b1011000001100011;
            15'b000001001101010 : data = 16'b1011000001110110;
            15'b000001001101011 : data = 16'b1011000010001001;
            15'b000001001101100 : data = 16'b1011000010011100;
            15'b000001001101101 : data = 16'b1011000010101111;
            15'b000001001101110 : data = 16'b1011000011000010;
            15'b000001001101111 : data = 16'b1011000011010101;
            15'b000001001110000 : data = 16'b1011000011101000;
            15'b000001001110001 : data = 16'b1011000011111011;
            15'b000001001110010 : data = 16'b1011000100001110;
            15'b000001001110011 : data = 16'b1011000100100001;
            15'b000001001110100 : data = 16'b1011000100110100;
            15'b000001001110101 : data = 16'b1011000101000111;
            15'b000001001110110 : data = 16'b1011000101011010;
            15'b000001001110111 : data = 16'b1011000101101101;
            15'b000001001111000 : data = 16'b1011000110000000;
            15'b000001001111001 : data = 16'b1011000110010011;
            15'b000001001111010 : data = 16'b1011000110100110;
            15'b000001001111011 : data = 16'b1011000110111001;
            15'b000001001111100 : data = 16'b1011000111001100;
            15'b000001001111101 : data = 16'b1011000111011111;
            15'b000001001111110 : data = 16'b1011000111110010;
            15'b000001001111111 : data = 16'b1011001000000101;
            15'b000001010000000 : data = 16'b1011001000011000;
            15'b000001010000001 : data = 16'b1011001000101011;
            15'b000001010000010 : data = 16'b1011001000111110;
            15'b000001010000011 : data = 16'b1011001001010000;
            15'b000001010000100 : data = 16'b1011001001100011;
            15'b000001010000101 : data = 16'b1011001001110110;
            15'b000001010000110 : data = 16'b1011001010001001;
            15'b000001010000111 : data = 16'b1011001010011100;
            15'b000001010001000 : data = 16'b1011001010101111;
            15'b000001010001001 : data = 16'b1011001011000010;
            15'b000001010001010 : data = 16'b1011001011010101;
            15'b000001010001011 : data = 16'b1011001011101000;
            15'b000001010001100 : data = 16'b1011001011111011;
            15'b000001010001101 : data = 16'b1011001100001110;
            15'b000001010001110 : data = 16'b1011001100100000;
            15'b000001010001111 : data = 16'b1011001100110011;
            15'b000001010010000 : data = 16'b1011001101000110;
            15'b000001010010001 : data = 16'b1011001101011001;
            15'b000001010010010 : data = 16'b1011001101101100;
            15'b000001010010011 : data = 16'b1011001101111111;
            15'b000001010010100 : data = 16'b1011001110010010;
            15'b000001010010101 : data = 16'b1011001110100100;
            15'b000001010010110 : data = 16'b1011001110110111;
            15'b000001010010111 : data = 16'b1011001111001010;
            15'b000001010011000 : data = 16'b1011001111011101;
            15'b000001010011001 : data = 16'b1011001111110000;
            15'b000001010011010 : data = 16'b1011010000000010;
            15'b000001010011011 : data = 16'b1011010000010101;
            15'b000001010011100 : data = 16'b1011010000101000;
            15'b000001010011101 : data = 16'b1011010000111011;
            15'b000001010011110 : data = 16'b1011010001001110;
            15'b000001010011111 : data = 16'b1011010001100000;
            15'b000001010100000 : data = 16'b1011010001110011;
            15'b000001010100001 : data = 16'b1011010010000110;
            15'b000001010100010 : data = 16'b1011010010011001;
            15'b000001010100011 : data = 16'b1011010010101100;
            15'b000001010100100 : data = 16'b1011010010111110;
            15'b000001010100101 : data = 16'b1011010011010001;
            15'b000001010100110 : data = 16'b1011010011100100;
            15'b000001010100111 : data = 16'b1011010011110111;
            15'b000001010101000 : data = 16'b1011010100001001;
            15'b000001010101001 : data = 16'b1011010100011100;
            15'b000001010101010 : data = 16'b1011010100101111;
            15'b000001010101011 : data = 16'b1011010101000010;
            15'b000001010101100 : data = 16'b1011010101010100;
            15'b000001010101101 : data = 16'b1011010101100111;
            15'b000001010101110 : data = 16'b1011010101111010;
            15'b000001010101111 : data = 16'b1011010110001100;
            15'b000001010110000 : data = 16'b1011010110011111;
            15'b000001010110001 : data = 16'b1011010110110010;
            15'b000001010110010 : data = 16'b1011010111000100;
            15'b000001010110011 : data = 16'b1011010111010111;
            15'b000001010110100 : data = 16'b1011010111101010;
            15'b000001010110101 : data = 16'b1011010111111100;
            15'b000001010110110 : data = 16'b1011011000001111;
            15'b000001010110111 : data = 16'b1011011000100010;
            15'b000001010111000 : data = 16'b1011011000110100;
            15'b000001010111001 : data = 16'b1011011001000111;
            15'b000001010111010 : data = 16'b1011011001011010;
            15'b000001010111011 : data = 16'b1011011001101100;
            15'b000001010111100 : data = 16'b1011011001111111;
            15'b000001010111101 : data = 16'b1011011010010010;
            15'b000001010111110 : data = 16'b1011011010100100;
            15'b000001010111111 : data = 16'b1011011010110111;
            15'b000001011000000 : data = 16'b1011011011001001;
            15'b000001011000001 : data = 16'b1011011011011100;
            15'b000001011000010 : data = 16'b1011011011101111;
            15'b000001011000011 : data = 16'b1011011100000001;
            15'b000001011000100 : data = 16'b1011011100010100;
            15'b000001011000101 : data = 16'b1011011100100110;
            15'b000001011000110 : data = 16'b1011011100111001;
            15'b000001011000111 : data = 16'b1011011101001100;
            15'b000001011001000 : data = 16'b1011011101011110;
            15'b000001011001001 : data = 16'b1011011101110001;
            15'b000001011001010 : data = 16'b1011011110000011;
            15'b000001011001011 : data = 16'b1011011110010110;
            15'b000001011001100 : data = 16'b1011011110101000;
            15'b000001011001101 : data = 16'b1011011110111011;
            15'b000001011001110 : data = 16'b1011011111001101;
            15'b000001011001111 : data = 16'b1011011111100000;
            15'b000001011010000 : data = 16'b1011011111110010;
            15'b000001011010001 : data = 16'b1011100000000101;
            15'b000001011010010 : data = 16'b1011100000010111;
            15'b000001011010011 : data = 16'b1011100000101010;
            15'b000001011010100 : data = 16'b1011100000111100;
            15'b000001011010101 : data = 16'b1011100001001111;
            15'b000001011010110 : data = 16'b1011100001100001;
            15'b000001011010111 : data = 16'b1011100001110100;
            15'b000001011011000 : data = 16'b1011100010000110;
            15'b000001011011001 : data = 16'b1011100010011001;
            15'b000001011011010 : data = 16'b1011100010101011;
            15'b000001011011011 : data = 16'b1011100010111110;
            15'b000001011011100 : data = 16'b1011100011010000;
            15'b000001011011101 : data = 16'b1011100011100011;
            15'b000001011011110 : data = 16'b1011100011110101;
            15'b000001011011111 : data = 16'b1011100100001000;
            15'b000001011100000 : data = 16'b1011100100011010;
            15'b000001011100001 : data = 16'b1011100100101100;
            15'b000001011100010 : data = 16'b1011100100111111;
            15'b000001011100011 : data = 16'b1011100101010001;
            15'b000001011100100 : data = 16'b1011100101100100;
            15'b000001011100101 : data = 16'b1011100101110110;
            15'b000001011100110 : data = 16'b1011100110001000;
            15'b000001011100111 : data = 16'b1011100110011011;
            15'b000001011101000 : data = 16'b1011100110101101;
            15'b000001011101001 : data = 16'b1011100111000000;
            15'b000001011101010 : data = 16'b1011100111010010;
            15'b000001011101011 : data = 16'b1011100111100100;
            15'b000001011101100 : data = 16'b1011100111110111;
            15'b000001011101101 : data = 16'b1011101000001001;
            15'b000001011101110 : data = 16'b1011101000011011;
            15'b000001011101111 : data = 16'b1011101000101110;
            15'b000001011110000 : data = 16'b1011101001000000;
            15'b000001011110001 : data = 16'b1011101001010010;
            15'b000001011110010 : data = 16'b1011101001100101;
            15'b000001011110011 : data = 16'b1011101001110111;
            15'b000001011110100 : data = 16'b1011101010001001;
            15'b000001011110101 : data = 16'b1011101010011100;
            15'b000001011110110 : data = 16'b1011101010101110;
            15'b000001011110111 : data = 16'b1011101011000000;
            15'b000001011111000 : data = 16'b1011101011010011;
            15'b000001011111001 : data = 16'b1011101011100101;
            15'b000001011111010 : data = 16'b1011101011110111;
            15'b000001011111011 : data = 16'b1011101100001001;
            15'b000001011111100 : data = 16'b1011101100011100;
            15'b000001011111101 : data = 16'b1011101100101110;
            15'b000001011111110 : data = 16'b1011101101000000;
            15'b000001011111111 : data = 16'b1011101101010010;
            15'b000001100000000 : data = 16'b1011101101100101;
            15'b000001100000001 : data = 16'b1011101101110111;
            15'b000001100000010 : data = 16'b1011101110001001;
            15'b000001100000011 : data = 16'b1011101110011011;
            15'b000001100000100 : data = 16'b1011101110101110;
            15'b000001100000101 : data = 16'b1011101111000000;
            15'b000001100000110 : data = 16'b1011101111010010;
            15'b000001100000111 : data = 16'b1011101111100100;
            15'b000001100001000 : data = 16'b1011101111110110;
            15'b000001100001001 : data = 16'b1011110000001001;
            15'b000001100001010 : data = 16'b1011110000011011;
            15'b000001100001011 : data = 16'b1011110000101101;
            15'b000001100001100 : data = 16'b1011110000111111;
            15'b000001100001101 : data = 16'b1011110001010001;
            15'b000001100001110 : data = 16'b1011110001100011;
            15'b000001100001111 : data = 16'b1011110001110110;
            15'b000001100010000 : data = 16'b1011110010001000;
            15'b000001100010001 : data = 16'b1011110010011010;
            15'b000001100010010 : data = 16'b1011110010101100;
            15'b000001100010011 : data = 16'b1011110010111110;
            15'b000001100010100 : data = 16'b1011110011010000;
            15'b000001100010101 : data = 16'b1011110011100010;
            15'b000001100010110 : data = 16'b1011110011110100;
            15'b000001100010111 : data = 16'b1011110100000110;
            15'b000001100011000 : data = 16'b1011110100011001;
            15'b000001100011001 : data = 16'b1011110100101011;
            15'b000001100011010 : data = 16'b1011110100111101;
            15'b000001100011011 : data = 16'b1011110101001111;
            15'b000001100011100 : data = 16'b1011110101100001;
            15'b000001100011101 : data = 16'b1011110101110011;
            15'b000001100011110 : data = 16'b1011110110000101;
            15'b000001100011111 : data = 16'b1011110110010111;
            15'b000001100100000 : data = 16'b1011110110101001;
            15'b000001100100001 : data = 16'b1011110110111011;
            15'b000001100100010 : data = 16'b1011110111001101;
            15'b000001100100011 : data = 16'b1011110111011111;
            15'b000001100100100 : data = 16'b1011110111110001;
            15'b000001100100101 : data = 16'b1011111000000011;
            15'b000001100100110 : data = 16'b1011111000010101;
            15'b000001100100111 : data = 16'b1011111000100111;
            15'b000001100101000 : data = 16'b1011111000111001;
            15'b000001100101001 : data = 16'b1011111001001011;
            15'b000001100101010 : data = 16'b1011111001011101;
            15'b000001100101011 : data = 16'b1011111001101111;
            15'b000001100101100 : data = 16'b1011111010000001;
            15'b000001100101101 : data = 16'b1011111010010011;
            15'b000001100101110 : data = 16'b1011111010100101;
            15'b000001100101111 : data = 16'b1011111010110111;
            15'b000001100110000 : data = 16'b1011111011001001;
            15'b000001100110001 : data = 16'b1011111011011011;
            15'b000001100110010 : data = 16'b1011111011101101;
            15'b000001100110011 : data = 16'b1011111011111111;
            15'b000001100110100 : data = 16'b1011111100010001;
            15'b000001100110101 : data = 16'b1011111100100011;
            15'b000001100110110 : data = 16'b1011111100110101;
            15'b000001100110111 : data = 16'b1011111101000110;
            15'b000001100111000 : data = 16'b1011111101011000;
            15'b000001100111001 : data = 16'b1011111101101010;
            15'b000001100111010 : data = 16'b1011111101111100;
            15'b000001100111011 : data = 16'b1011111110001110;
            15'b000001100111100 : data = 16'b1011111110100000;
            15'b000001100111101 : data = 16'b1011111110110010;
            15'b000001100111110 : data = 16'b1011111111000100;
            15'b000001100111111 : data = 16'b1011111111010101;
            15'b000001101000000 : data = 16'b1011111111100111;
            15'b000001101000001 : data = 16'b1011111111111001;
            15'b000001101000010 : data = 16'b1100000000001011;
            15'b000001101000011 : data = 16'b1100000000011101;
            15'b000001101000100 : data = 16'b1100000000101111;
            15'b000001101000101 : data = 16'b1100000001000000;
            15'b000001101000110 : data = 16'b1100000001010010;
            15'b000001101000111 : data = 16'b1100000001100100;
            15'b000001101001000 : data = 16'b1100000001110110;
            15'b000001101001001 : data = 16'b1100000010001000;
            15'b000001101001010 : data = 16'b1100000010011001;
            15'b000001101001011 : data = 16'b1100000010101011;
            15'b000001101001100 : data = 16'b1100000010111101;
            15'b000001101001101 : data = 16'b1100000011001111;
            15'b000001101001110 : data = 16'b1100000011100000;
            15'b000001101001111 : data = 16'b1100000011110010;
            15'b000001101010000 : data = 16'b1100000100000100;
            15'b000001101010001 : data = 16'b1100000100010110;
            15'b000001101010010 : data = 16'b1100000100100111;
            15'b000001101010011 : data = 16'b1100000100111001;
            15'b000001101010100 : data = 16'b1100000101001011;
            15'b000001101010101 : data = 16'b1100000101011100;
            15'b000001101010110 : data = 16'b1100000101101110;
            15'b000001101010111 : data = 16'b1100000110000000;
            15'b000001101011000 : data = 16'b1100000110010001;
            15'b000001101011001 : data = 16'b1100000110100011;
            15'b000001101011010 : data = 16'b1100000110110101;
            15'b000001101011011 : data = 16'b1100000111000110;
            15'b000001101011100 : data = 16'b1100000111011000;
            15'b000001101011101 : data = 16'b1100000111101010;
            15'b000001101011110 : data = 16'b1100000111111011;
            15'b000001101011111 : data = 16'b1100001000001101;
            15'b000001101100000 : data = 16'b1100001000011111;
            15'b000001101100001 : data = 16'b1100001000110000;
            15'b000001101100010 : data = 16'b1100001001000010;
            15'b000001101100011 : data = 16'b1100001001010100;
            15'b000001101100100 : data = 16'b1100001001100101;
            15'b000001101100101 : data = 16'b1100001001110111;
            15'b000001101100110 : data = 16'b1100001010001000;
            15'b000001101100111 : data = 16'b1100001010011010;
            15'b000001101101000 : data = 16'b1100001010101100;
            15'b000001101101001 : data = 16'b1100001010111101;
            15'b000001101101010 : data = 16'b1100001011001111;
            15'b000001101101011 : data = 16'b1100001011100000;
            15'b000001101101100 : data = 16'b1100001011110010;
            15'b000001101101101 : data = 16'b1100001100000011;
            15'b000001101101110 : data = 16'b1100001100010101;
            15'b000001101101111 : data = 16'b1100001100100110;
            15'b000001101110000 : data = 16'b1100001100111000;
            15'b000001101110001 : data = 16'b1100001101001001;
            15'b000001101110010 : data = 16'b1100001101011011;
            15'b000001101110011 : data = 16'b1100001101101100;
            15'b000001101110100 : data = 16'b1100001101111110;
            15'b000001101110101 : data = 16'b1100001110001111;
            15'b000001101110110 : data = 16'b1100001110100001;
            15'b000001101110111 : data = 16'b1100001110110010;
            15'b000001101111000 : data = 16'b1100001111000100;
            15'b000001101111001 : data = 16'b1100001111010101;
            15'b000001101111010 : data = 16'b1100001111100111;
            15'b000001101111011 : data = 16'b1100001111111000;
            15'b000001101111100 : data = 16'b1100010000001010;
            15'b000001101111101 : data = 16'b1100010000011011;
            15'b000001101111110 : data = 16'b1100010000101101;
            15'b000001101111111 : data = 16'b1100010000111110;
            15'b000001110000000 : data = 16'b1100010001001111;
            15'b000001110000001 : data = 16'b1100010001100001;
            15'b000001110000010 : data = 16'b1100010001110010;
            15'b000001110000011 : data = 16'b1100010010000100;
            15'b000001110000100 : data = 16'b1100010010010101;
            15'b000001110000101 : data = 16'b1100010010100110;
            15'b000001110000110 : data = 16'b1100010010111000;
            15'b000001110000111 : data = 16'b1100010011001001;
            15'b000001110001000 : data = 16'b1100010011011010;
            15'b000001110001001 : data = 16'b1100010011101100;
            15'b000001110001010 : data = 16'b1100010011111101;
            15'b000001110001011 : data = 16'b1100010100001110;
            15'b000001110001100 : data = 16'b1100010100100000;
            15'b000001110001101 : data = 16'b1100010100110001;
            15'b000001110001110 : data = 16'b1100010101000010;
            15'b000001110001111 : data = 16'b1100010101010100;
            15'b000001110010000 : data = 16'b1100010101100101;
            15'b000001110010001 : data = 16'b1100010101110110;
            15'b000001110010010 : data = 16'b1100010110001000;
            15'b000001110010011 : data = 16'b1100010110011001;
            15'b000001110010100 : data = 16'b1100010110101010;
            15'b000001110010101 : data = 16'b1100010110111011;
            15'b000001110010110 : data = 16'b1100010111001101;
            15'b000001110010111 : data = 16'b1100010111011110;
            15'b000001110011000 : data = 16'b1100010111101111;
            15'b000001110011001 : data = 16'b1100011000000000;
            15'b000001110011010 : data = 16'b1100011000010010;
            15'b000001110011011 : data = 16'b1100011000100011;
            15'b000001110011100 : data = 16'b1100011000110100;
            15'b000001110011101 : data = 16'b1100011001000101;
            15'b000001110011110 : data = 16'b1100011001010111;
            15'b000001110011111 : data = 16'b1100011001101000;
            15'b000001110100000 : data = 16'b1100011001111001;
            15'b000001110100001 : data = 16'b1100011010001010;
            15'b000001110100010 : data = 16'b1100011010011011;
            15'b000001110100011 : data = 16'b1100011010101100;
            15'b000001110100100 : data = 16'b1100011010111110;
            15'b000001110100101 : data = 16'b1100011011001111;
            15'b000001110100110 : data = 16'b1100011011100000;
            15'b000001110100111 : data = 16'b1100011011110001;
            15'b000001110101000 : data = 16'b1100011100000010;
            15'b000001110101001 : data = 16'b1100011100010011;
            15'b000001110101010 : data = 16'b1100011100100100;
            15'b000001110101011 : data = 16'b1100011100110110;
            15'b000001110101100 : data = 16'b1100011101000111;
            15'b000001110101101 : data = 16'b1100011101011000;
            15'b000001110101110 : data = 16'b1100011101101001;
            15'b000001110101111 : data = 16'b1100011101111010;
            15'b000001110110000 : data = 16'b1100011110001011;
            15'b000001110110001 : data = 16'b1100011110011100;
            15'b000001110110010 : data = 16'b1100011110101101;
            15'b000001110110011 : data = 16'b1100011110111110;
            15'b000001110110100 : data = 16'b1100011111001111;
            15'b000001110110101 : data = 16'b1100011111100000;
            15'b000001110110110 : data = 16'b1100011111110001;
            15'b000001110110111 : data = 16'b1100100000000010;
            15'b000001110111000 : data = 16'b1100100000010011;
            15'b000001110111001 : data = 16'b1100100000100100;
            15'b000001110111010 : data = 16'b1100100000110101;
            15'b000001110111011 : data = 16'b1100100001000110;
            15'b000001110111100 : data = 16'b1100100001010111;
            15'b000001110111101 : data = 16'b1100100001101000;
            15'b000001110111110 : data = 16'b1100100001111001;
            15'b000001110111111 : data = 16'b1100100010001010;
            15'b000001111000000 : data = 16'b1100100010011011;
            15'b000001111000001 : data = 16'b1100100010101100;
            15'b000001111000010 : data = 16'b1100100010111101;
            15'b000001111000011 : data = 16'b1100100011001110;
            15'b000001111000100 : data = 16'b1100100011011111;
            15'b000001111000101 : data = 16'b1100100011110000;
            15'b000001111000110 : data = 16'b1100100100000001;
            15'b000001111000111 : data = 16'b1100100100010010;
            15'b000001111001000 : data = 16'b1100100100100011;
            15'b000001111001001 : data = 16'b1100100100110011;
            15'b000001111001010 : data = 16'b1100100101000100;
            15'b000001111001011 : data = 16'b1100100101010101;
            15'b000001111001100 : data = 16'b1100100101100110;
            15'b000001111001101 : data = 16'b1100100101110111;
            15'b000001111001110 : data = 16'b1100100110001000;
            15'b000001111001111 : data = 16'b1100100110011001;
            15'b000001111010000 : data = 16'b1100100110101010;
            15'b000001111010001 : data = 16'b1100100110111010;
            15'b000001111010010 : data = 16'b1100100111001011;
            15'b000001111010011 : data = 16'b1100100111011100;
            15'b000001111010100 : data = 16'b1100100111101101;
            15'b000001111010101 : data = 16'b1100100111111110;
            15'b000001111010110 : data = 16'b1100101000001110;
            15'b000001111010111 : data = 16'b1100101000011111;
            15'b000001111011000 : data = 16'b1100101000110000;
            15'b000001111011001 : data = 16'b1100101001000001;
            15'b000001111011010 : data = 16'b1100101001010010;
            15'b000001111011011 : data = 16'b1100101001100010;
            15'b000001111011100 : data = 16'b1100101001110011;
            15'b000001111011101 : data = 16'b1100101010000100;
            15'b000001111011110 : data = 16'b1100101010010101;
            15'b000001111011111 : data = 16'b1100101010100101;
            15'b000001111100000 : data = 16'b1100101010110110;
            15'b000001111100001 : data = 16'b1100101011000111;
            15'b000001111100010 : data = 16'b1100101011010111;
            15'b000001111100011 : data = 16'b1100101011101000;
            15'b000001111100100 : data = 16'b1100101011111001;
            15'b000001111100101 : data = 16'b1100101100001001;
            15'b000001111100110 : data = 16'b1100101100011010;
            15'b000001111100111 : data = 16'b1100101100101011;
            15'b000001111101000 : data = 16'b1100101100111011;
            15'b000001111101001 : data = 16'b1100101101001100;
            15'b000001111101010 : data = 16'b1100101101011101;
            15'b000001111101011 : data = 16'b1100101101101101;
            15'b000001111101100 : data = 16'b1100101101111110;
            15'b000001111101101 : data = 16'b1100101110001111;
            15'b000001111101110 : data = 16'b1100101110011111;
            15'b000001111101111 : data = 16'b1100101110110000;
            15'b000001111110000 : data = 16'b1100101111000000;
            15'b000001111110001 : data = 16'b1100101111010001;
            15'b000001111110010 : data = 16'b1100101111100010;
            15'b000001111110011 : data = 16'b1100101111110010;
            15'b000001111110100 : data = 16'b1100110000000011;
            15'b000001111110101 : data = 16'b1100110000010011;
            15'b000001111110110 : data = 16'b1100110000100100;
            15'b000001111110111 : data = 16'b1100110000110100;
            15'b000001111111000 : data = 16'b1100110001000101;
            15'b000001111111001 : data = 16'b1100110001010110;
            15'b000001111111010 : data = 16'b1100110001100110;
            15'b000001111111011 : data = 16'b1100110001110111;
            15'b000001111111100 : data = 16'b1100110010000111;
            15'b000001111111101 : data = 16'b1100110010011000;
            15'b000001111111110 : data = 16'b1100110010101000;
            15'b000001111111111 : data = 16'b1100110010111001;
            15'b000010000000000 : data = 16'b1100110011001001;
            15'b000010000000001 : data = 16'b1100110011011001;
            15'b000010000000010 : data = 16'b1100110011101010;
            15'b000010000000011 : data = 16'b1100110011111010;
            15'b000010000000100 : data = 16'b1100110100001011;
            15'b000010000000101 : data = 16'b1100110100011011;
            15'b000010000000110 : data = 16'b1100110100101100;
            15'b000010000000111 : data = 16'b1100110100111100;
            15'b000010000001000 : data = 16'b1100110101001101;
            15'b000010000001001 : data = 16'b1100110101011101;
            15'b000010000001010 : data = 16'b1100110101101101;
            15'b000010000001011 : data = 16'b1100110101111110;
            15'b000010000001100 : data = 16'b1100110110001110;
            15'b000010000001101 : data = 16'b1100110110011110;
            15'b000010000001110 : data = 16'b1100110110101111;
            15'b000010000001111 : data = 16'b1100110110111111;
            15'b000010000010000 : data = 16'b1100110111010000;
            15'b000010000010001 : data = 16'b1100110111100000;
            15'b000010000010010 : data = 16'b1100110111110000;
            15'b000010000010011 : data = 16'b1100111000000001;
            15'b000010000010100 : data = 16'b1100111000010001;
            15'b000010000010101 : data = 16'b1100111000100001;
            15'b000010000010110 : data = 16'b1100111000110001;
            15'b000010000010111 : data = 16'b1100111001000010;
            15'b000010000011000 : data = 16'b1100111001010010;
            15'b000010000011001 : data = 16'b1100111001100010;
            15'b000010000011010 : data = 16'b1100111001110011;
            15'b000010000011011 : data = 16'b1100111010000011;
            15'b000010000011100 : data = 16'b1100111010010011;
            15'b000010000011101 : data = 16'b1100111010100011;
            15'b000010000011110 : data = 16'b1100111010110100;
            15'b000010000011111 : data = 16'b1100111011000100;
            15'b000010000100000 : data = 16'b1100111011010100;
            15'b000010000100001 : data = 16'b1100111011100100;
            15'b000010000100010 : data = 16'b1100111011110101;
            15'b000010000100011 : data = 16'b1100111100000101;
            15'b000010000100100 : data = 16'b1100111100010101;
            15'b000010000100101 : data = 16'b1100111100100101;
            15'b000010000100110 : data = 16'b1100111100110101;
            15'b000010000100111 : data = 16'b1100111101000101;
            15'b000010000101000 : data = 16'b1100111101010110;
            15'b000010000101001 : data = 16'b1100111101100110;
            15'b000010000101010 : data = 16'b1100111101110110;
            15'b000010000101011 : data = 16'b1100111110000110;
            15'b000010000101100 : data = 16'b1100111110010110;
            15'b000010000101101 : data = 16'b1100111110100110;
            15'b000010000101110 : data = 16'b1100111110110110;
            15'b000010000101111 : data = 16'b1100111111000110;
            15'b000010000110000 : data = 16'b1100111111010111;
            15'b000010000110001 : data = 16'b1100111111100111;
            15'b000010000110010 : data = 16'b1100111111110111;
            15'b000010000110011 : data = 16'b1101000000000111;
            15'b000010000110100 : data = 16'b1101000000010111;
            15'b000010000110101 : data = 16'b1101000000100111;
            15'b000010000110110 : data = 16'b1101000000110111;
            15'b000010000110111 : data = 16'b1101000001000111;
            15'b000010000111000 : data = 16'b1101000001010111;
            15'b000010000111001 : data = 16'b1101000001100111;
            15'b000010000111010 : data = 16'b1101000001110111;
            15'b000010000111011 : data = 16'b1101000010000111;
            15'b000010000111100 : data = 16'b1101000010010111;
            15'b000010000111101 : data = 16'b1101000010100111;
            15'b000010000111110 : data = 16'b1101000010110111;
            15'b000010000111111 : data = 16'b1101000011000111;
            15'b000010001000000 : data = 16'b1101000011010111;
            15'b000010001000001 : data = 16'b1101000011100111;
            15'b000010001000010 : data = 16'b1101000011110111;
            15'b000010001000011 : data = 16'b1101000100000111;
            15'b000010001000100 : data = 16'b1101000100010111;
            15'b000010001000101 : data = 16'b1101000100100111;
            15'b000010001000110 : data = 16'b1101000100110111;
            15'b000010001000111 : data = 16'b1101000101000111;
            15'b000010001001000 : data = 16'b1101000101010110;
            15'b000010001001001 : data = 16'b1101000101100110;
            15'b000010001001010 : data = 16'b1101000101110110;
            15'b000010001001011 : data = 16'b1101000110000110;
            15'b000010001001100 : data = 16'b1101000110010110;
            15'b000010001001101 : data = 16'b1101000110100110;
            15'b000010001001110 : data = 16'b1101000110110110;
            15'b000010001001111 : data = 16'b1101000111000110;
            15'b000010001010000 : data = 16'b1101000111010101;
            15'b000010001010001 : data = 16'b1101000111100101;
            15'b000010001010010 : data = 16'b1101000111110101;
            15'b000010001010011 : data = 16'b1101001000000101;
            15'b000010001010100 : data = 16'b1101001000010101;
            15'b000010001010101 : data = 16'b1101001000100100;
            15'b000010001010110 : data = 16'b1101001000110100;
            15'b000010001010111 : data = 16'b1101001001000100;
            15'b000010001011000 : data = 16'b1101001001010100;
            15'b000010001011001 : data = 16'b1101001001100011;
            15'b000010001011010 : data = 16'b1101001001110011;
            15'b000010001011011 : data = 16'b1101001010000011;
            15'b000010001011100 : data = 16'b1101001010010011;
            15'b000010001011101 : data = 16'b1101001010100010;
            15'b000010001011110 : data = 16'b1101001010110010;
            15'b000010001011111 : data = 16'b1101001011000010;
            15'b000010001100000 : data = 16'b1101001011010010;
            15'b000010001100001 : data = 16'b1101001011100001;
            15'b000010001100010 : data = 16'b1101001011110001;
            15'b000010001100011 : data = 16'b1101001100000001;
            15'b000010001100100 : data = 16'b1101001100010000;
            15'b000010001100101 : data = 16'b1101001100100000;
            15'b000010001100110 : data = 16'b1101001100110000;
            15'b000010001100111 : data = 16'b1101001100111111;
            15'b000010001101000 : data = 16'b1101001101001111;
            15'b000010001101001 : data = 16'b1101001101011111;
            15'b000010001101010 : data = 16'b1101001101101110;
            15'b000010001101011 : data = 16'b1101001101111110;
            15'b000010001101100 : data = 16'b1101001110001101;
            15'b000010001101101 : data = 16'b1101001110011101;
            15'b000010001101110 : data = 16'b1101001110101101;
            15'b000010001101111 : data = 16'b1101001110111100;
            15'b000010001110000 : data = 16'b1101001111001100;
            15'b000010001110001 : data = 16'b1101001111011011;
            15'b000010001110010 : data = 16'b1101001111101011;
            15'b000010001110011 : data = 16'b1101001111111010;
            15'b000010001110100 : data = 16'b1101010000001010;
            15'b000010001110101 : data = 16'b1101010000011001;
            15'b000010001110110 : data = 16'b1101010000101001;
            15'b000010001110111 : data = 16'b1101010000111000;
            15'b000010001111000 : data = 16'b1101010001001000;
            15'b000010001111001 : data = 16'b1101010001010111;
            15'b000010001111010 : data = 16'b1101010001100111;
            15'b000010001111011 : data = 16'b1101010001110110;
            15'b000010001111100 : data = 16'b1101010010000110;
            15'b000010001111101 : data = 16'b1101010010010101;
            15'b000010001111110 : data = 16'b1101010010100101;
            15'b000010001111111 : data = 16'b1101010010110100;
            15'b000010010000000 : data = 16'b1101010011000100;
            15'b000010010000001 : data = 16'b1101010011010011;
            15'b000010010000010 : data = 16'b1101010011100010;
            15'b000010010000011 : data = 16'b1101010011110010;
            15'b000010010000100 : data = 16'b1101010100000001;
            15'b000010010000101 : data = 16'b1101010100010001;
            15'b000010010000110 : data = 16'b1101010100100000;
            15'b000010010000111 : data = 16'b1101010100101111;
            15'b000010010001000 : data = 16'b1101010100111111;
            15'b000010010001001 : data = 16'b1101010101001110;
            15'b000010010001010 : data = 16'b1101010101011101;
            15'b000010010001011 : data = 16'b1101010101101101;
            15'b000010010001100 : data = 16'b1101010101111100;
            15'b000010010001101 : data = 16'b1101010110001011;
            15'b000010010001110 : data = 16'b1101010110011011;
            15'b000010010001111 : data = 16'b1101010110101010;
            15'b000010010010000 : data = 16'b1101010110111001;
            15'b000010010010001 : data = 16'b1101010111001001;
            15'b000010010010010 : data = 16'b1101010111011000;
            15'b000010010010011 : data = 16'b1101010111100111;
            15'b000010010010100 : data = 16'b1101010111110110;
            15'b000010010010101 : data = 16'b1101011000000110;
            15'b000010010010110 : data = 16'b1101011000010101;
            15'b000010010010111 : data = 16'b1101011000100100;
            15'b000010010011000 : data = 16'b1101011000110011;
            15'b000010010011001 : data = 16'b1101011001000011;
            15'b000010010011010 : data = 16'b1101011001010010;
            15'b000010010011011 : data = 16'b1101011001100001;
            15'b000010010011100 : data = 16'b1101011001110000;
            15'b000010010011101 : data = 16'b1101011001111111;
            15'b000010010011110 : data = 16'b1101011010001110;
            15'b000010010011111 : data = 16'b1101011010011110;
            15'b000010010100000 : data = 16'b1101011010101101;
            15'b000010010100001 : data = 16'b1101011010111100;
            15'b000010010100010 : data = 16'b1101011011001011;
            15'b000010010100011 : data = 16'b1101011011011010;
            15'b000010010100100 : data = 16'b1101011011101001;
            15'b000010010100101 : data = 16'b1101011011111000;
            15'b000010010100110 : data = 16'b1101011100001000;
            15'b000010010100111 : data = 16'b1101011100010111;
            15'b000010010101000 : data = 16'b1101011100100110;
            15'b000010010101001 : data = 16'b1101011100110101;
            15'b000010010101010 : data = 16'b1101011101000100;
            15'b000010010101011 : data = 16'b1101011101010011;
            15'b000010010101100 : data = 16'b1101011101100010;
            15'b000010010101101 : data = 16'b1101011101110001;
            15'b000010010101110 : data = 16'b1101011110000000;
            15'b000010010101111 : data = 16'b1101011110001111;
            15'b000010010110000 : data = 16'b1101011110011110;
            15'b000010010110001 : data = 16'b1101011110101101;
            15'b000010010110010 : data = 16'b1101011110111100;
            15'b000010010110011 : data = 16'b1101011111001011;
            15'b000010010110100 : data = 16'b1101011111011010;
            15'b000010010110101 : data = 16'b1101011111101001;
            15'b000010010110110 : data = 16'b1101011111111000;
            15'b000010010110111 : data = 16'b1101100000000111;
            15'b000010010111000 : data = 16'b1101100000010110;
            15'b000010010111001 : data = 16'b1101100000100101;
            15'b000010010111010 : data = 16'b1101100000110100;
            15'b000010010111011 : data = 16'b1101100001000011;
            15'b000010010111100 : data = 16'b1101100001010010;
            15'b000010010111101 : data = 16'b1101100001100000;
            15'b000010010111110 : data = 16'b1101100001101111;
            15'b000010010111111 : data = 16'b1101100001111110;
            15'b000010011000000 : data = 16'b1101100010001101;
            15'b000010011000001 : data = 16'b1101100010011100;
            15'b000010011000010 : data = 16'b1101100010101011;
            15'b000010011000011 : data = 16'b1101100010111010;
            15'b000010011000100 : data = 16'b1101100011001000;
            15'b000010011000101 : data = 16'b1101100011010111;
            15'b000010011000110 : data = 16'b1101100011100110;
            15'b000010011000111 : data = 16'b1101100011110101;
            15'b000010011001000 : data = 16'b1101100100000100;
            15'b000010011001001 : data = 16'b1101100100010010;
            15'b000010011001010 : data = 16'b1101100100100001;
            15'b000010011001011 : data = 16'b1101100100110000;
            15'b000010011001100 : data = 16'b1101100100111111;
            15'b000010011001101 : data = 16'b1101100101001110;
            15'b000010011001110 : data = 16'b1101100101011100;
            15'b000010011001111 : data = 16'b1101100101101011;
            15'b000010011010000 : data = 16'b1101100101111010;
            15'b000010011010001 : data = 16'b1101100110001000;
            15'b000010011010010 : data = 16'b1101100110010111;
            15'b000010011010011 : data = 16'b1101100110100110;
            15'b000010011010100 : data = 16'b1101100110110101;
            15'b000010011010101 : data = 16'b1101100111000011;
            15'b000010011010110 : data = 16'b1101100111010010;
            15'b000010011010111 : data = 16'b1101100111100001;
            15'b000010011011000 : data = 16'b1101100111101111;
            15'b000010011011001 : data = 16'b1101100111111110;
            15'b000010011011010 : data = 16'b1101101000001101;
            15'b000010011011011 : data = 16'b1101101000011011;
            15'b000010011011100 : data = 16'b1101101000101010;
            15'b000010011011101 : data = 16'b1101101000111000;
            15'b000010011011110 : data = 16'b1101101001000111;
            15'b000010011011111 : data = 16'b1101101001010110;
            15'b000010011100000 : data = 16'b1101101001100100;
            15'b000010011100001 : data = 16'b1101101001110011;
            15'b000010011100010 : data = 16'b1101101010000001;
            15'b000010011100011 : data = 16'b1101101010010000;
            15'b000010011100100 : data = 16'b1101101010011110;
            15'b000010011100101 : data = 16'b1101101010101101;
            15'b000010011100110 : data = 16'b1101101010111011;
            15'b000010011100111 : data = 16'b1101101011001010;
            15'b000010011101000 : data = 16'b1101101011011000;
            15'b000010011101001 : data = 16'b1101101011100111;
            15'b000010011101010 : data = 16'b1101101011110101;
            15'b000010011101011 : data = 16'b1101101100000100;
            15'b000010011101100 : data = 16'b1101101100010010;
            15'b000010011101101 : data = 16'b1101101100100001;
            15'b000010011101110 : data = 16'b1101101100101111;
            15'b000010011101111 : data = 16'b1101101100111110;
            15'b000010011110000 : data = 16'b1101101101001100;
            15'b000010011110001 : data = 16'b1101101101011011;
            15'b000010011110010 : data = 16'b1101101101101001;
            15'b000010011110011 : data = 16'b1101101101110111;
            15'b000010011110100 : data = 16'b1101101110000110;
            15'b000010011110101 : data = 16'b1101101110010100;
            15'b000010011110110 : data = 16'b1101101110100011;
            15'b000010011110111 : data = 16'b1101101110110001;
            15'b000010011111000 : data = 16'b1101101110111111;
            15'b000010011111001 : data = 16'b1101101111001110;
            15'b000010011111010 : data = 16'b1101101111011100;
            15'b000010011111011 : data = 16'b1101101111101010;
            15'b000010011111100 : data = 16'b1101101111111001;
            15'b000010011111101 : data = 16'b1101110000000111;
            15'b000010011111110 : data = 16'b1101110000010101;
            15'b000010011111111 : data = 16'b1101110000100100;
            15'b000010100000000 : data = 16'b1101110000110010;
            15'b000010100000001 : data = 16'b1101110001000000;
            15'b000010100000010 : data = 16'b1101110001001110;
            15'b000010100000011 : data = 16'b1101110001011101;
            15'b000010100000100 : data = 16'b1101110001101011;
            15'b000010100000101 : data = 16'b1101110001111001;
            15'b000010100000110 : data = 16'b1101110010000111;
            15'b000010100000111 : data = 16'b1101110010010110;
            15'b000010100001000 : data = 16'b1101110010100100;
            15'b000010100001001 : data = 16'b1101110010110010;
            15'b000010100001010 : data = 16'b1101110011000000;
            15'b000010100001011 : data = 16'b1101110011001110;
            15'b000010100001100 : data = 16'b1101110011011101;
            15'b000010100001101 : data = 16'b1101110011101011;
            15'b000010100001110 : data = 16'b1101110011111001;
            15'b000010100001111 : data = 16'b1101110100000111;
            15'b000010100010000 : data = 16'b1101110100010101;
            15'b000010100010001 : data = 16'b1101110100100011;
            15'b000010100010010 : data = 16'b1101110100110001;
            15'b000010100010011 : data = 16'b1101110101000000;
            15'b000010100010100 : data = 16'b1101110101001110;
            15'b000010100010101 : data = 16'b1101110101011100;
            15'b000010100010110 : data = 16'b1101110101101010;
            15'b000010100010111 : data = 16'b1101110101111000;
            15'b000010100011000 : data = 16'b1101110110000110;
            15'b000010100011001 : data = 16'b1101110110010100;
            15'b000010100011010 : data = 16'b1101110110100010;
            15'b000010100011011 : data = 16'b1101110110110000;
            15'b000010100011100 : data = 16'b1101110110111110;
            15'b000010100011101 : data = 16'b1101110111001100;
            15'b000010100011110 : data = 16'b1101110111011010;
            15'b000010100011111 : data = 16'b1101110111101000;
            15'b000010100100000 : data = 16'b1101110111110110;
            15'b000010100100001 : data = 16'b1101111000000100;
            15'b000010100100010 : data = 16'b1101111000010010;
            15'b000010100100011 : data = 16'b1101111000100000;
            15'b000010100100100 : data = 16'b1101111000101110;
            15'b000010100100101 : data = 16'b1101111000111100;
            15'b000010100100110 : data = 16'b1101111001001010;
            15'b000010100100111 : data = 16'b1101111001011000;
            15'b000010100101000 : data = 16'b1101111001100110;
            15'b000010100101001 : data = 16'b1101111001110011;
            15'b000010100101010 : data = 16'b1101111010000001;
            15'b000010100101011 : data = 16'b1101111010001111;
            15'b000010100101100 : data = 16'b1101111010011101;
            15'b000010100101101 : data = 16'b1101111010101011;
            15'b000010100101110 : data = 16'b1101111010111001;
            15'b000010100101111 : data = 16'b1101111011000111;
            15'b000010100110000 : data = 16'b1101111011010101;
            15'b000010100110001 : data = 16'b1101111011100010;
            15'b000010100110010 : data = 16'b1101111011110000;
            15'b000010100110011 : data = 16'b1101111011111110;
            15'b000010100110100 : data = 16'b1101111100001100;
            15'b000010100110101 : data = 16'b1101111100011010;
            15'b000010100110110 : data = 16'b1101111100100111;
            15'b000010100110111 : data = 16'b1101111100110101;
            15'b000010100111000 : data = 16'b1101111101000011;
            15'b000010100111001 : data = 16'b1101111101010001;
            15'b000010100111010 : data = 16'b1101111101011110;
            15'b000010100111011 : data = 16'b1101111101101100;
            15'b000010100111100 : data = 16'b1101111101111010;
            15'b000010100111101 : data = 16'b1101111110000111;
            15'b000010100111110 : data = 16'b1101111110010101;
            15'b000010100111111 : data = 16'b1101111110100011;
            15'b000010101000000 : data = 16'b1101111110110001;
            15'b000010101000001 : data = 16'b1101111110111110;
            15'b000010101000010 : data = 16'b1101111111001100;
            15'b000010101000011 : data = 16'b1101111111011010;
            15'b000010101000100 : data = 16'b1101111111100111;
            15'b000010101000101 : data = 16'b1101111111110101;
            15'b000010101000110 : data = 16'b1110000000000010;
            15'b000010101000111 : data = 16'b1110000000010000;
            15'b000010101001000 : data = 16'b1110000000011110;
            15'b000010101001001 : data = 16'b1110000000101011;
            15'b000010101001010 : data = 16'b1110000000111001;
            15'b000010101001011 : data = 16'b1110000001000110;
            15'b000010101001100 : data = 16'b1110000001010100;
            15'b000010101001101 : data = 16'b1110000001100001;
            15'b000010101001110 : data = 16'b1110000001101111;
            15'b000010101001111 : data = 16'b1110000001111101;
            15'b000010101010000 : data = 16'b1110000010001010;
            15'b000010101010001 : data = 16'b1110000010011000;
            15'b000010101010010 : data = 16'b1110000010100101;
            15'b000010101010011 : data = 16'b1110000010110011;
            15'b000010101010100 : data = 16'b1110000011000000;
            15'b000010101010101 : data = 16'b1110000011001110;
            15'b000010101010110 : data = 16'b1110000011011011;
            15'b000010101010111 : data = 16'b1110000011101000;
            15'b000010101011000 : data = 16'b1110000011110110;
            15'b000010101011001 : data = 16'b1110000100000011;
            15'b000010101011010 : data = 16'b1110000100010001;
            15'b000010101011011 : data = 16'b1110000100011110;
            15'b000010101011100 : data = 16'b1110000100101100;
            15'b000010101011101 : data = 16'b1110000100111001;
            15'b000010101011110 : data = 16'b1110000101000110;
            15'b000010101011111 : data = 16'b1110000101010100;
            15'b000010101100000 : data = 16'b1110000101100001;
            15'b000010101100001 : data = 16'b1110000101101110;
            15'b000010101100010 : data = 16'b1110000101111100;
            15'b000010101100011 : data = 16'b1110000110001001;
            15'b000010101100100 : data = 16'b1110000110010110;
            15'b000010101100101 : data = 16'b1110000110100100;
            15'b000010101100110 : data = 16'b1110000110110001;
            15'b000010101100111 : data = 16'b1110000110111110;
            15'b000010101101000 : data = 16'b1110000111001100;
            15'b000010101101001 : data = 16'b1110000111011001;
            15'b000010101101010 : data = 16'b1110000111100110;
            15'b000010101101011 : data = 16'b1110000111110011;
            15'b000010101101100 : data = 16'b1110001000000001;
            15'b000010101101101 : data = 16'b1110001000001110;
            15'b000010101101110 : data = 16'b1110001000011011;
            15'b000010101101111 : data = 16'b1110001000101000;
            15'b000010101110000 : data = 16'b1110001000110110;
            15'b000010101110001 : data = 16'b1110001001000011;
            15'b000010101110010 : data = 16'b1110001001010000;
            15'b000010101110011 : data = 16'b1110001001011101;
            15'b000010101110100 : data = 16'b1110001001101010;
            15'b000010101110101 : data = 16'b1110001001110111;
            15'b000010101110110 : data = 16'b1110001010000101;
            15'b000010101110111 : data = 16'b1110001010010010;
            15'b000010101111000 : data = 16'b1110001010011111;
            15'b000010101111001 : data = 16'b1110001010101100;
            15'b000010101111010 : data = 16'b1110001010111001;
            15'b000010101111011 : data = 16'b1110001011000110;
            15'b000010101111100 : data = 16'b1110001011010011;
            15'b000010101111101 : data = 16'b1110001011100000;
            15'b000010101111110 : data = 16'b1110001011101101;
            15'b000010101111111 : data = 16'b1110001011111011;
            15'b000010110000000 : data = 16'b1110001100001000;
            15'b000010110000001 : data = 16'b1110001100010101;
            15'b000010110000010 : data = 16'b1110001100100010;
            15'b000010110000011 : data = 16'b1110001100101111;
            15'b000010110000100 : data = 16'b1110001100111100;
            15'b000010110000101 : data = 16'b1110001101001001;
            15'b000010110000110 : data = 16'b1110001101010110;
            15'b000010110000111 : data = 16'b1110001101100011;
            15'b000010110001000 : data = 16'b1110001101110000;
            15'b000010110001001 : data = 16'b1110001101111101;
            15'b000010110001010 : data = 16'b1110001110001010;
            15'b000010110001011 : data = 16'b1110001110010110;
            15'b000010110001100 : data = 16'b1110001110100011;
            15'b000010110001101 : data = 16'b1110001110110000;
            15'b000010110001110 : data = 16'b1110001110111101;
            15'b000010110001111 : data = 16'b1110001111001010;
            15'b000010110010000 : data = 16'b1110001111010111;
            15'b000010110010001 : data = 16'b1110001111100100;
            15'b000010110010010 : data = 16'b1110001111110001;
            15'b000010110010011 : data = 16'b1110001111111110;
            15'b000010110010100 : data = 16'b1110010000001010;
            15'b000010110010101 : data = 16'b1110010000010111;
            15'b000010110010110 : data = 16'b1110010000100100;
            15'b000010110010111 : data = 16'b1110010000110001;
            15'b000010110011000 : data = 16'b1110010000111110;
            15'b000010110011001 : data = 16'b1110010001001011;
            15'b000010110011010 : data = 16'b1110010001010111;
            15'b000010110011011 : data = 16'b1110010001100100;
            15'b000010110011100 : data = 16'b1110010001110001;
            15'b000010110011101 : data = 16'b1110010001111110;
            15'b000010110011110 : data = 16'b1110010010001010;
            15'b000010110011111 : data = 16'b1110010010010111;
            15'b000010110100000 : data = 16'b1110010010100100;
            15'b000010110100001 : data = 16'b1110010010110001;
            15'b000010110100010 : data = 16'b1110010010111101;
            15'b000010110100011 : data = 16'b1110010011001010;
            15'b000010110100100 : data = 16'b1110010011010111;
            15'b000010110100101 : data = 16'b1110010011100011;
            15'b000010110100110 : data = 16'b1110010011110000;
            15'b000010110100111 : data = 16'b1110010011111101;
            15'b000010110101000 : data = 16'b1110010100001001;
            15'b000010110101001 : data = 16'b1110010100010110;
            15'b000010110101010 : data = 16'b1110010100100011;
            15'b000010110101011 : data = 16'b1110010100101111;
            15'b000010110101100 : data = 16'b1110010100111100;
            15'b000010110101101 : data = 16'b1110010101001000;
            15'b000010110101110 : data = 16'b1110010101010101;
            15'b000010110101111 : data = 16'b1110010101100001;
            15'b000010110110000 : data = 16'b1110010101101110;
            15'b000010110110001 : data = 16'b1110010101111011;
            15'b000010110110010 : data = 16'b1110010110000111;
            15'b000010110110011 : data = 16'b1110010110010100;
            15'b000010110110100 : data = 16'b1110010110100000;
            15'b000010110110101 : data = 16'b1110010110101101;
            15'b000010110110110 : data = 16'b1110010110111001;
            15'b000010110110111 : data = 16'b1110010111000110;
            15'b000010110111000 : data = 16'b1110010111010010;
            15'b000010110111001 : data = 16'b1110010111011111;
            15'b000010110111010 : data = 16'b1110010111101011;
            15'b000010110111011 : data = 16'b1110010111111000;
            15'b000010110111100 : data = 16'b1110011000000100;
            15'b000010110111101 : data = 16'b1110011000010000;
            15'b000010110111110 : data = 16'b1110011000011101;
            15'b000010110111111 : data = 16'b1110011000101001;
            15'b000010111000000 : data = 16'b1110011000110110;
            15'b000010111000001 : data = 16'b1110011001000010;
            15'b000010111000010 : data = 16'b1110011001001110;
            15'b000010111000011 : data = 16'b1110011001011011;
            15'b000010111000100 : data = 16'b1110011001100111;
            15'b000010111000101 : data = 16'b1110011001110011;
            15'b000010111000110 : data = 16'b1110011010000000;
            15'b000010111000111 : data = 16'b1110011010001100;
            15'b000010111001000 : data = 16'b1110011010011000;
            15'b000010111001001 : data = 16'b1110011010100101;
            15'b000010111001010 : data = 16'b1110011010110001;
            15'b000010111001011 : data = 16'b1110011010111101;
            15'b000010111001100 : data = 16'b1110011011001010;
            15'b000010111001101 : data = 16'b1110011011010110;
            15'b000010111001110 : data = 16'b1110011011100010;
            15'b000010111001111 : data = 16'b1110011011101110;
            15'b000010111010000 : data = 16'b1110011011111011;
            15'b000010111010001 : data = 16'b1110011100000111;
            15'b000010111010010 : data = 16'b1110011100010011;
            15'b000010111010011 : data = 16'b1110011100011111;
            15'b000010111010100 : data = 16'b1110011100101011;
            15'b000010111010101 : data = 16'b1110011100111000;
            15'b000010111010110 : data = 16'b1110011101000100;
            15'b000010111010111 : data = 16'b1110011101010000;
            15'b000010111011000 : data = 16'b1110011101011100;
            15'b000010111011001 : data = 16'b1110011101101000;
            15'b000010111011010 : data = 16'b1110011101110100;
            15'b000010111011011 : data = 16'b1110011110000000;
            15'b000010111011100 : data = 16'b1110011110001101;
            15'b000010111011101 : data = 16'b1110011110011001;
            15'b000010111011110 : data = 16'b1110011110100101;
            15'b000010111011111 : data = 16'b1110011110110001;
            15'b000010111100000 : data = 16'b1110011110111101;
            15'b000010111100001 : data = 16'b1110011111001001;
            15'b000010111100010 : data = 16'b1110011111010101;
            15'b000010111100011 : data = 16'b1110011111100001;
            15'b000010111100100 : data = 16'b1110011111101101;
            15'b000010111100101 : data = 16'b1110011111111001;
            15'b000010111100110 : data = 16'b1110100000000101;
            15'b000010111100111 : data = 16'b1110100000010001;
            15'b000010111101000 : data = 16'b1110100000011101;
            15'b000010111101001 : data = 16'b1110100000101001;
            15'b000010111101010 : data = 16'b1110100000110101;
            15'b000010111101011 : data = 16'b1110100001000001;
            15'b000010111101100 : data = 16'b1110100001001101;
            15'b000010111101101 : data = 16'b1110100001011001;
            15'b000010111101110 : data = 16'b1110100001100101;
            15'b000010111101111 : data = 16'b1110100001110001;
            15'b000010111110000 : data = 16'b1110100001111100;
            15'b000010111110001 : data = 16'b1110100010001000;
            15'b000010111110010 : data = 16'b1110100010010100;
            15'b000010111110011 : data = 16'b1110100010100000;
            15'b000010111110100 : data = 16'b1110100010101100;
            15'b000010111110101 : data = 16'b1110100010111000;
            15'b000010111110110 : data = 16'b1110100011000100;
            15'b000010111110111 : data = 16'b1110100011001111;
            15'b000010111111000 : data = 16'b1110100011011011;
            15'b000010111111001 : data = 16'b1110100011100111;
            15'b000010111111010 : data = 16'b1110100011110011;
            15'b000010111111011 : data = 16'b1110100011111111;
            15'b000010111111100 : data = 16'b1110100100001010;
            15'b000010111111101 : data = 16'b1110100100010110;
            15'b000010111111110 : data = 16'b1110100100100010;
            15'b000010111111111 : data = 16'b1110100100101110;
            15'b000011000000000 : data = 16'b1110100100111001;
            15'b000011000000001 : data = 16'b1110100101000101;
            15'b000011000000010 : data = 16'b1110100101010001;
            15'b000011000000011 : data = 16'b1110100101011101;
            15'b000011000000100 : data = 16'b1110100101101000;
            15'b000011000000101 : data = 16'b1110100101110100;
            15'b000011000000110 : data = 16'b1110100110000000;
            15'b000011000000111 : data = 16'b1110100110001011;
            15'b000011000001000 : data = 16'b1110100110010111;
            15'b000011000001001 : data = 16'b1110100110100010;
            15'b000011000001010 : data = 16'b1110100110101110;
            15'b000011000001011 : data = 16'b1110100110111010;
            15'b000011000001100 : data = 16'b1110100111000101;
            15'b000011000001101 : data = 16'b1110100111010001;
            15'b000011000001110 : data = 16'b1110100111011100;
            15'b000011000001111 : data = 16'b1110100111101000;
            15'b000011000010000 : data = 16'b1110100111110100;
            15'b000011000010001 : data = 16'b1110100111111111;
            15'b000011000010010 : data = 16'b1110101000001011;
            15'b000011000010011 : data = 16'b1110101000010110;
            15'b000011000010100 : data = 16'b1110101000100010;
            15'b000011000010101 : data = 16'b1110101000101101;
            15'b000011000010110 : data = 16'b1110101000111001;
            15'b000011000010111 : data = 16'b1110101001000100;
            15'b000011000011000 : data = 16'b1110101001010000;
            15'b000011000011001 : data = 16'b1110101001011011;
            15'b000011000011010 : data = 16'b1110101001100111;
            15'b000011000011011 : data = 16'b1110101001110010;
            15'b000011000011100 : data = 16'b1110101001111101;
            15'b000011000011101 : data = 16'b1110101010001001;
            15'b000011000011110 : data = 16'b1110101010010100;
            15'b000011000011111 : data = 16'b1110101010100000;
            15'b000011000100000 : data = 16'b1110101010101011;
            15'b000011000100001 : data = 16'b1110101010110110;
            15'b000011000100010 : data = 16'b1110101011000010;
            15'b000011000100011 : data = 16'b1110101011001101;
            15'b000011000100100 : data = 16'b1110101011011000;
            15'b000011000100101 : data = 16'b1110101011100100;
            15'b000011000100110 : data = 16'b1110101011101111;
            15'b000011000100111 : data = 16'b1110101011111010;
            15'b000011000101000 : data = 16'b1110101100000110;
            15'b000011000101001 : data = 16'b1110101100010001;
            15'b000011000101010 : data = 16'b1110101100011100;
            15'b000011000101011 : data = 16'b1110101100101000;
            15'b000011000101100 : data = 16'b1110101100110011;
            15'b000011000101101 : data = 16'b1110101100111110;
            15'b000011000101110 : data = 16'b1110101101001001;
            15'b000011000101111 : data = 16'b1110101101010100;
            15'b000011000110000 : data = 16'b1110101101100000;
            15'b000011000110001 : data = 16'b1110101101101011;
            15'b000011000110010 : data = 16'b1110101101110110;
            15'b000011000110011 : data = 16'b1110101110000001;
            15'b000011000110100 : data = 16'b1110101110001100;
            15'b000011000110101 : data = 16'b1110101110011000;
            15'b000011000110110 : data = 16'b1110101110100011;
            15'b000011000110111 : data = 16'b1110101110101110;
            15'b000011000111000 : data = 16'b1110101110111001;
            15'b000011000111001 : data = 16'b1110101111000100;
            15'b000011000111010 : data = 16'b1110101111001111;
            15'b000011000111011 : data = 16'b1110101111011010;
            15'b000011000111100 : data = 16'b1110101111100101;
            15'b000011000111101 : data = 16'b1110101111110000;
            15'b000011000111110 : data = 16'b1110101111111100;
            15'b000011000111111 : data = 16'b1110110000000111;
            15'b000011001000000 : data = 16'b1110110000010010;
            15'b000011001000001 : data = 16'b1110110000011101;
            15'b000011001000010 : data = 16'b1110110000101000;
            15'b000011001000011 : data = 16'b1110110000110011;
            15'b000011001000100 : data = 16'b1110110000111110;
            15'b000011001000101 : data = 16'b1110110001001001;
            15'b000011001000110 : data = 16'b1110110001010100;
            15'b000011001000111 : data = 16'b1110110001011111;
            15'b000011001001000 : data = 16'b1110110001101001;
            15'b000011001001001 : data = 16'b1110110001110100;
            15'b000011001001010 : data = 16'b1110110001111111;
            15'b000011001001011 : data = 16'b1110110010001010;
            15'b000011001001100 : data = 16'b1110110010010101;
            15'b000011001001101 : data = 16'b1110110010100000;
            15'b000011001001110 : data = 16'b1110110010101011;
            15'b000011001001111 : data = 16'b1110110010110110;
            15'b000011001010000 : data = 16'b1110110011000001;
            15'b000011001010001 : data = 16'b1110110011001100;
            15'b000011001010010 : data = 16'b1110110011010110;
            15'b000011001010011 : data = 16'b1110110011100001;
            15'b000011001010100 : data = 16'b1110110011101100;
            15'b000011001010101 : data = 16'b1110110011110111;
            15'b000011001010110 : data = 16'b1110110100000010;
            15'b000011001010111 : data = 16'b1110110100001100;
            15'b000011001011000 : data = 16'b1110110100010111;
            15'b000011001011001 : data = 16'b1110110100100010;
            15'b000011001011010 : data = 16'b1110110100101101;
            15'b000011001011011 : data = 16'b1110110100110111;
            15'b000011001011100 : data = 16'b1110110101000010;
            15'b000011001011101 : data = 16'b1110110101001101;
            15'b000011001011110 : data = 16'b1110110101011000;
            15'b000011001011111 : data = 16'b1110110101100010;
            15'b000011001100000 : data = 16'b1110110101101101;
            15'b000011001100001 : data = 16'b1110110101111000;
            15'b000011001100010 : data = 16'b1110110110000010;
            15'b000011001100011 : data = 16'b1110110110001101;
            15'b000011001100100 : data = 16'b1110110110011000;
            15'b000011001100101 : data = 16'b1110110110100010;
            15'b000011001100110 : data = 16'b1110110110101101;
            15'b000011001100111 : data = 16'b1110110110110111;
            15'b000011001101000 : data = 16'b1110110111000010;
            15'b000011001101001 : data = 16'b1110110111001101;
            15'b000011001101010 : data = 16'b1110110111010111;
            15'b000011001101011 : data = 16'b1110110111100010;
            15'b000011001101100 : data = 16'b1110110111101100;
            15'b000011001101101 : data = 16'b1110110111110111;
            15'b000011001101110 : data = 16'b1110111000000001;
            15'b000011001101111 : data = 16'b1110111000001100;
            15'b000011001110000 : data = 16'b1110111000010110;
            15'b000011001110001 : data = 16'b1110111000100001;
            15'b000011001110010 : data = 16'b1110111000101011;
            15'b000011001110011 : data = 16'b1110111000110110;
            15'b000011001110100 : data = 16'b1110111001000000;
            15'b000011001110101 : data = 16'b1110111001001011;
            15'b000011001110110 : data = 16'b1110111001010101;
            15'b000011001110111 : data = 16'b1110111001100000;
            15'b000011001111000 : data = 16'b1110111001101010;
            15'b000011001111001 : data = 16'b1110111001110101;
            15'b000011001111010 : data = 16'b1110111001111111;
            15'b000011001111011 : data = 16'b1110111010001001;
            15'b000011001111100 : data = 16'b1110111010010100;
            15'b000011001111101 : data = 16'b1110111010011110;
            15'b000011001111110 : data = 16'b1110111010101000;
            15'b000011001111111 : data = 16'b1110111010110011;
            15'b000011010000000 : data = 16'b1110111010111101;
            15'b000011010000001 : data = 16'b1110111011000111;
            15'b000011010000010 : data = 16'b1110111011010010;
            15'b000011010000011 : data = 16'b1110111011011100;
            15'b000011010000100 : data = 16'b1110111011100110;
            15'b000011010000101 : data = 16'b1110111011110001;
            15'b000011010000110 : data = 16'b1110111011111011;
            15'b000011010000111 : data = 16'b1110111100000101;
            15'b000011010001000 : data = 16'b1110111100001111;
            15'b000011010001001 : data = 16'b1110111100011010;
            15'b000011010001010 : data = 16'b1110111100100100;
            15'b000011010001011 : data = 16'b1110111100101110;
            15'b000011010001100 : data = 16'b1110111100111000;
            15'b000011010001101 : data = 16'b1110111101000010;
            15'b000011010001110 : data = 16'b1110111101001100;
            15'b000011010001111 : data = 16'b1110111101010111;
            15'b000011010010000 : data = 16'b1110111101100001;
            15'b000011010010001 : data = 16'b1110111101101011;
            15'b000011010010010 : data = 16'b1110111101110101;
            15'b000011010010011 : data = 16'b1110111101111111;
            15'b000011010010100 : data = 16'b1110111110001001;
            15'b000011010010101 : data = 16'b1110111110010011;
            15'b000011010010110 : data = 16'b1110111110011101;
            15'b000011010010111 : data = 16'b1110111110101000;
            15'b000011010011000 : data = 16'b1110111110110010;
            15'b000011010011001 : data = 16'b1110111110111100;
            15'b000011010011010 : data = 16'b1110111111000110;
            15'b000011010011011 : data = 16'b1110111111010000;
            15'b000011010011100 : data = 16'b1110111111011010;
            15'b000011010011101 : data = 16'b1110111111100100;
            15'b000011010011110 : data = 16'b1110111111101110;
            15'b000011010011111 : data = 16'b1110111111111000;
            15'b000011010100000 : data = 16'b1111000000000010;
            15'b000011010100001 : data = 16'b1111000000001100;
            15'b000011010100010 : data = 16'b1111000000010110;
            15'b000011010100011 : data = 16'b1111000000100000;
            15'b000011010100100 : data = 16'b1111000000101001;
            15'b000011010100101 : data = 16'b1111000000110011;
            15'b000011010100110 : data = 16'b1111000000111101;
            15'b000011010100111 : data = 16'b1111000001000111;
            15'b000011010101000 : data = 16'b1111000001010001;
            15'b000011010101001 : data = 16'b1111000001011011;
            15'b000011010101010 : data = 16'b1111000001100101;
            15'b000011010101011 : data = 16'b1111000001101111;
            15'b000011010101100 : data = 16'b1111000001111000;
            15'b000011010101101 : data = 16'b1111000010000010;
            15'b000011010101110 : data = 16'b1111000010001100;
            15'b000011010101111 : data = 16'b1111000010010110;
            15'b000011010110000 : data = 16'b1111000010100000;
            15'b000011010110001 : data = 16'b1111000010101001;
            15'b000011010110010 : data = 16'b1111000010110011;
            15'b000011010110011 : data = 16'b1111000010111101;
            15'b000011010110100 : data = 16'b1111000011000111;
            15'b000011010110101 : data = 16'b1111000011010000;
            15'b000011010110110 : data = 16'b1111000011011010;
            15'b000011010110111 : data = 16'b1111000011100100;
            15'b000011010111000 : data = 16'b1111000011101110;
            15'b000011010111001 : data = 16'b1111000011110111;
            15'b000011010111010 : data = 16'b1111000100000001;
            15'b000011010111011 : data = 16'b1111000100001011;
            15'b000011010111100 : data = 16'b1111000100010100;
            15'b000011010111101 : data = 16'b1111000100011110;
            15'b000011010111110 : data = 16'b1111000100100111;
            15'b000011010111111 : data = 16'b1111000100110001;
            15'b000011011000000 : data = 16'b1111000100111011;
            15'b000011011000001 : data = 16'b1111000101000100;
            15'b000011011000010 : data = 16'b1111000101001110;
            15'b000011011000011 : data = 16'b1111000101010111;
            15'b000011011000100 : data = 16'b1111000101100001;
            15'b000011011000101 : data = 16'b1111000101101011;
            15'b000011011000110 : data = 16'b1111000101110100;
            15'b000011011000111 : data = 16'b1111000101111110;
            15'b000011011001000 : data = 16'b1111000110000111;
            15'b000011011001001 : data = 16'b1111000110010001;
            15'b000011011001010 : data = 16'b1111000110011010;
            15'b000011011001011 : data = 16'b1111000110100100;
            15'b000011011001100 : data = 16'b1111000110101101;
            15'b000011011001101 : data = 16'b1111000110110111;
            15'b000011011001110 : data = 16'b1111000111000000;
            15'b000011011001111 : data = 16'b1111000111001001;
            15'b000011011010000 : data = 16'b1111000111010011;
            15'b000011011010001 : data = 16'b1111000111011100;
            15'b000011011010010 : data = 16'b1111000111100110;
            15'b000011011010011 : data = 16'b1111000111101111;
            15'b000011011010100 : data = 16'b1111000111111000;
            15'b000011011010101 : data = 16'b1111001000000010;
            15'b000011011010110 : data = 16'b1111001000001011;
            15'b000011011010111 : data = 16'b1111001000010100;
            15'b000011011011000 : data = 16'b1111001000011110;
            15'b000011011011001 : data = 16'b1111001000100111;
            15'b000011011011010 : data = 16'b1111001000110000;
            15'b000011011011011 : data = 16'b1111001000111010;
            15'b000011011011100 : data = 16'b1111001001000011;
            15'b000011011011101 : data = 16'b1111001001001100;
            15'b000011011011110 : data = 16'b1111001001010110;
            15'b000011011011111 : data = 16'b1111001001011111;
            15'b000011011100000 : data = 16'b1111001001101000;
            15'b000011011100001 : data = 16'b1111001001110001;
            15'b000011011100010 : data = 16'b1111001001111010;
            15'b000011011100011 : data = 16'b1111001010000100;
            15'b000011011100100 : data = 16'b1111001010001101;
            15'b000011011100101 : data = 16'b1111001010010110;
            15'b000011011100110 : data = 16'b1111001010011111;
            15'b000011011100111 : data = 16'b1111001010101000;
            15'b000011011101000 : data = 16'b1111001010110001;
            15'b000011011101001 : data = 16'b1111001010111011;
            15'b000011011101010 : data = 16'b1111001011000100;
            15'b000011011101011 : data = 16'b1111001011001101;
            15'b000011011101100 : data = 16'b1111001011010110;
            15'b000011011101101 : data = 16'b1111001011011111;
            15'b000011011101110 : data = 16'b1111001011101000;
            15'b000011011101111 : data = 16'b1111001011110001;
            15'b000011011110000 : data = 16'b1111001011111010;
            15'b000011011110001 : data = 16'b1111001100000011;
            15'b000011011110010 : data = 16'b1111001100001100;
            15'b000011011110011 : data = 16'b1111001100010101;
            15'b000011011110100 : data = 16'b1111001100011110;
            15'b000011011110101 : data = 16'b1111001100100111;
            15'b000011011110110 : data = 16'b1111001100110000;
            15'b000011011110111 : data = 16'b1111001100111001;
            15'b000011011111000 : data = 16'b1111001101000010;
            15'b000011011111001 : data = 16'b1111001101001011;
            15'b000011011111010 : data = 16'b1111001101010100;
            15'b000011011111011 : data = 16'b1111001101011101;
            15'b000011011111100 : data = 16'b1111001101100110;
            15'b000011011111101 : data = 16'b1111001101101111;
            15'b000011011111110 : data = 16'b1111001101111000;
            15'b000011011111111 : data = 16'b1111001110000001;
            15'b000011100000000 : data = 16'b1111001110001001;
            15'b000011100000001 : data = 16'b1111001110010010;
            15'b000011100000010 : data = 16'b1111001110011011;
            15'b000011100000011 : data = 16'b1111001110100100;
            15'b000011100000100 : data = 16'b1111001110101101;
            15'b000011100000101 : data = 16'b1111001110110110;
            15'b000011100000110 : data = 16'b1111001110111110;
            15'b000011100000111 : data = 16'b1111001111000111;
            15'b000011100001000 : data = 16'b1111001111010000;
            15'b000011100001001 : data = 16'b1111001111011001;
            15'b000011100001010 : data = 16'b1111001111100001;
            15'b000011100001011 : data = 16'b1111001111101010;
            15'b000011100001100 : data = 16'b1111001111110011;
            15'b000011100001101 : data = 16'b1111001111111100;
            15'b000011100001110 : data = 16'b1111010000000100;
            15'b000011100001111 : data = 16'b1111010000001101;
            15'b000011100010000 : data = 16'b1111010000010110;
            15'b000011100010001 : data = 16'b1111010000011110;
            15'b000011100010010 : data = 16'b1111010000100111;
            15'b000011100010011 : data = 16'b1111010000110000;
            15'b000011100010100 : data = 16'b1111010000111000;
            15'b000011100010101 : data = 16'b1111010001000001;
            15'b000011100010110 : data = 16'b1111010001001010;
            15'b000011100010111 : data = 16'b1111010001010010;
            15'b000011100011000 : data = 16'b1111010001011011;
            15'b000011100011001 : data = 16'b1111010001100011;
            15'b000011100011010 : data = 16'b1111010001101100;
            15'b000011100011011 : data = 16'b1111010001110100;
            15'b000011100011100 : data = 16'b1111010001111101;
            15'b000011100011101 : data = 16'b1111010010000101;
            15'b000011100011110 : data = 16'b1111010010001110;
            15'b000011100011111 : data = 16'b1111010010010110;
            15'b000011100100000 : data = 16'b1111010010011111;
            15'b000011100100001 : data = 16'b1111010010100111;
            15'b000011100100010 : data = 16'b1111010010110000;
            15'b000011100100011 : data = 16'b1111010010111000;
            15'b000011100100100 : data = 16'b1111010011000001;
            15'b000011100100101 : data = 16'b1111010011001001;
            15'b000011100100110 : data = 16'b1111010011010010;
            15'b000011100100111 : data = 16'b1111010011011010;
            15'b000011100101000 : data = 16'b1111010011100010;
            15'b000011100101001 : data = 16'b1111010011101011;
            15'b000011100101010 : data = 16'b1111010011110011;
            15'b000011100101011 : data = 16'b1111010011111100;
            15'b000011100101100 : data = 16'b1111010100000100;
            15'b000011100101101 : data = 16'b1111010100001100;
            15'b000011100101110 : data = 16'b1111010100010101;
            15'b000011100101111 : data = 16'b1111010100011101;
            15'b000011100110000 : data = 16'b1111010100100101;
            15'b000011100110001 : data = 16'b1111010100101101;
            15'b000011100110010 : data = 16'b1111010100110110;
            15'b000011100110011 : data = 16'b1111010100111110;
            15'b000011100110100 : data = 16'b1111010101000110;
            15'b000011100110101 : data = 16'b1111010101001111;
            15'b000011100110110 : data = 16'b1111010101010111;
            15'b000011100110111 : data = 16'b1111010101011111;
            15'b000011100111000 : data = 16'b1111010101100111;
            15'b000011100111001 : data = 16'b1111010101101111;
            15'b000011100111010 : data = 16'b1111010101111000;
            15'b000011100111011 : data = 16'b1111010110000000;
            15'b000011100111100 : data = 16'b1111010110001000;
            15'b000011100111101 : data = 16'b1111010110010000;
            15'b000011100111110 : data = 16'b1111010110011000;
            15'b000011100111111 : data = 16'b1111010110100000;
            15'b000011101000000 : data = 16'b1111010110101000;
            15'b000011101000001 : data = 16'b1111010110110001;
            15'b000011101000010 : data = 16'b1111010110111001;
            15'b000011101000011 : data = 16'b1111010111000001;
            15'b000011101000100 : data = 16'b1111010111001001;
            15'b000011101000101 : data = 16'b1111010111010001;
            15'b000011101000110 : data = 16'b1111010111011001;
            15'b000011101000111 : data = 16'b1111010111100001;
            15'b000011101001000 : data = 16'b1111010111101001;
            15'b000011101001001 : data = 16'b1111010111110001;
            15'b000011101001010 : data = 16'b1111010111111001;
            15'b000011101001011 : data = 16'b1111011000000001;
            15'b000011101001100 : data = 16'b1111011000001001;
            15'b000011101001101 : data = 16'b1111011000010001;
            15'b000011101001110 : data = 16'b1111011000011001;
            15'b000011101001111 : data = 16'b1111011000100001;
            15'b000011101010000 : data = 16'b1111011000101001;
            15'b000011101010001 : data = 16'b1111011000110000;
            15'b000011101010010 : data = 16'b1111011000111000;
            15'b000011101010011 : data = 16'b1111011001000000;
            15'b000011101010100 : data = 16'b1111011001001000;
            15'b000011101010101 : data = 16'b1111011001010000;
            15'b000011101010110 : data = 16'b1111011001011000;
            15'b000011101010111 : data = 16'b1111011001100000;
            15'b000011101011000 : data = 16'b1111011001101000;
            15'b000011101011001 : data = 16'b1111011001101111;
            15'b000011101011010 : data = 16'b1111011001110111;
            15'b000011101011011 : data = 16'b1111011001111111;
            15'b000011101011100 : data = 16'b1111011010000111;
            15'b000011101011101 : data = 16'b1111011010001110;
            15'b000011101011110 : data = 16'b1111011010010110;
            15'b000011101011111 : data = 16'b1111011010011110;
            15'b000011101100000 : data = 16'b1111011010100110;
            15'b000011101100001 : data = 16'b1111011010101101;
            15'b000011101100010 : data = 16'b1111011010110101;
            15'b000011101100011 : data = 16'b1111011010111101;
            15'b000011101100100 : data = 16'b1111011011000100;
            15'b000011101100101 : data = 16'b1111011011001100;
            15'b000011101100110 : data = 16'b1111011011010100;
            15'b000011101100111 : data = 16'b1111011011011011;
            15'b000011101101000 : data = 16'b1111011011100011;
            15'b000011101101001 : data = 16'b1111011011101011;
            15'b000011101101010 : data = 16'b1111011011110010;
            15'b000011101101011 : data = 16'b1111011011111010;
            15'b000011101101100 : data = 16'b1111011100000001;
            15'b000011101101101 : data = 16'b1111011100001001;
            15'b000011101101110 : data = 16'b1111011100010001;
            15'b000011101101111 : data = 16'b1111011100011000;
            15'b000011101110000 : data = 16'b1111011100100000;
            15'b000011101110001 : data = 16'b1111011100100111;
            15'b000011101110010 : data = 16'b1111011100101111;
            15'b000011101110011 : data = 16'b1111011100110110;
            15'b000011101110100 : data = 16'b1111011100111110;
            15'b000011101110101 : data = 16'b1111011101000101;
            15'b000011101110110 : data = 16'b1111011101001101;
            15'b000011101110111 : data = 16'b1111011101010100;
            15'b000011101111000 : data = 16'b1111011101011100;
            15'b000011101111001 : data = 16'b1111011101100011;
            15'b000011101111010 : data = 16'b1111011101101010;
            15'b000011101111011 : data = 16'b1111011101110010;
            15'b000011101111100 : data = 16'b1111011101111001;
            15'b000011101111101 : data = 16'b1111011110000001;
            15'b000011101111110 : data = 16'b1111011110001000;
            15'b000011101111111 : data = 16'b1111011110001111;
            15'b000011110000000 : data = 16'b1111011110010111;
            15'b000011110000001 : data = 16'b1111011110011110;
            15'b000011110000010 : data = 16'b1111011110100101;
            15'b000011110000011 : data = 16'b1111011110101101;
            15'b000011110000100 : data = 16'b1111011110110100;
            15'b000011110000101 : data = 16'b1111011110111011;
            15'b000011110000110 : data = 16'b1111011111000010;
            15'b000011110000111 : data = 16'b1111011111001010;
            15'b000011110001000 : data = 16'b1111011111010001;
            15'b000011110001001 : data = 16'b1111011111011000;
            15'b000011110001010 : data = 16'b1111011111011111;
            15'b000011110001011 : data = 16'b1111011111100111;
            15'b000011110001100 : data = 16'b1111011111101110;
            15'b000011110001101 : data = 16'b1111011111110101;
            15'b000011110001110 : data = 16'b1111011111111100;
            15'b000011110001111 : data = 16'b1111100000000011;
            15'b000011110010000 : data = 16'b1111100000001011;
            15'b000011110010001 : data = 16'b1111100000010010;
            15'b000011110010010 : data = 16'b1111100000011001;
            15'b000011110010011 : data = 16'b1111100000100000;
            15'b000011110010100 : data = 16'b1111100000100111;
            15'b000011110010101 : data = 16'b1111100000101110;
            15'b000011110010110 : data = 16'b1111100000110101;
            15'b000011110010111 : data = 16'b1111100000111100;
            15'b000011110011000 : data = 16'b1111100001000011;
            15'b000011110011001 : data = 16'b1111100001001010;
            15'b000011110011010 : data = 16'b1111100001010001;
            15'b000011110011011 : data = 16'b1111100001011000;
            15'b000011110011100 : data = 16'b1111100001011111;
            15'b000011110011101 : data = 16'b1111100001100110;
            15'b000011110011110 : data = 16'b1111100001101101;
            15'b000011110011111 : data = 16'b1111100001110100;
            15'b000011110100000 : data = 16'b1111100001111011;
            15'b000011110100001 : data = 16'b1111100010000010;
            15'b000011110100010 : data = 16'b1111100010001001;
            15'b000011110100011 : data = 16'b1111100010010000;
            15'b000011110100100 : data = 16'b1111100010010111;
            15'b000011110100101 : data = 16'b1111100010011110;
            15'b000011110100110 : data = 16'b1111100010100101;
            15'b000011110100111 : data = 16'b1111100010101100;
            15'b000011110101000 : data = 16'b1111100010110010;
            15'b000011110101001 : data = 16'b1111100010111001;
            15'b000011110101010 : data = 16'b1111100011000000;
            15'b000011110101011 : data = 16'b1111100011000111;
            15'b000011110101100 : data = 16'b1111100011001110;
            15'b000011110101101 : data = 16'b1111100011010101;
            15'b000011110101110 : data = 16'b1111100011011011;
            15'b000011110101111 : data = 16'b1111100011100010;
            15'b000011110110000 : data = 16'b1111100011101001;
            15'b000011110110001 : data = 16'b1111100011110000;
            15'b000011110110010 : data = 16'b1111100011110110;
            15'b000011110110011 : data = 16'b1111100011111101;
            15'b000011110110100 : data = 16'b1111100100000100;
            15'b000011110110101 : data = 16'b1111100100001011;
            15'b000011110110110 : data = 16'b1111100100010001;
            15'b000011110110111 : data = 16'b1111100100011000;
            15'b000011110111000 : data = 16'b1111100100011111;
            15'b000011110111001 : data = 16'b1111100100100101;
            15'b000011110111010 : data = 16'b1111100100101100;
            15'b000011110111011 : data = 16'b1111100100110010;
            15'b000011110111100 : data = 16'b1111100100111001;
            15'b000011110111101 : data = 16'b1111100101000000;
            15'b000011110111110 : data = 16'b1111100101000110;
            15'b000011110111111 : data = 16'b1111100101001101;
            15'b000011111000000 : data = 16'b1111100101010011;
            15'b000011111000001 : data = 16'b1111100101011010;
            15'b000011111000010 : data = 16'b1111100101100000;
            15'b000011111000011 : data = 16'b1111100101100111;
            15'b000011111000100 : data = 16'b1111100101101110;
            15'b000011111000101 : data = 16'b1111100101110100;
            15'b000011111000110 : data = 16'b1111100101111011;
            15'b000011111000111 : data = 16'b1111100110000001;
            15'b000011111001000 : data = 16'b1111100110000111;
            15'b000011111001001 : data = 16'b1111100110001110;
            15'b000011111001010 : data = 16'b1111100110010100;
            15'b000011111001011 : data = 16'b1111100110011011;
            15'b000011111001100 : data = 16'b1111100110100001;
            15'b000011111001101 : data = 16'b1111100110101000;
            15'b000011111001110 : data = 16'b1111100110101110;
            15'b000011111001111 : data = 16'b1111100110110100;
            15'b000011111010000 : data = 16'b1111100110111011;
            15'b000011111010001 : data = 16'b1111100111000001;
            15'b000011111010010 : data = 16'b1111100111000111;
            15'b000011111010011 : data = 16'b1111100111001110;
            15'b000011111010100 : data = 16'b1111100111010100;
            15'b000011111010101 : data = 16'b1111100111011010;
            15'b000011111010110 : data = 16'b1111100111100001;
            15'b000011111010111 : data = 16'b1111100111100111;
            15'b000011111011000 : data = 16'b1111100111101101;
            15'b000011111011001 : data = 16'b1111100111110100;
            15'b000011111011010 : data = 16'b1111100111111010;
            15'b000011111011011 : data = 16'b1111101000000000;
            15'b000011111011100 : data = 16'b1111101000000110;
            15'b000011111011101 : data = 16'b1111101000001100;
            15'b000011111011110 : data = 16'b1111101000010011;
            15'b000011111011111 : data = 16'b1111101000011001;
            15'b000011111100000 : data = 16'b1111101000011111;
            15'b000011111100001 : data = 16'b1111101000100101;
            15'b000011111100010 : data = 16'b1111101000101011;
            15'b000011111100011 : data = 16'b1111101000110001;
            15'b000011111100100 : data = 16'b1111101000111000;
            15'b000011111100101 : data = 16'b1111101000111110;
            15'b000011111100110 : data = 16'b1111101001000100;
            15'b000011111100111 : data = 16'b1111101001001010;
            15'b000011111101000 : data = 16'b1111101001010000;
            15'b000011111101001 : data = 16'b1111101001010110;
            15'b000011111101010 : data = 16'b1111101001011100;
            15'b000011111101011 : data = 16'b1111101001100010;
            15'b000011111101100 : data = 16'b1111101001101000;
            15'b000011111101101 : data = 16'b1111101001101110;
            15'b000011111101110 : data = 16'b1111101001110100;
            15'b000011111101111 : data = 16'b1111101001111010;
            15'b000011111110000 : data = 16'b1111101010000000;
            15'b000011111110001 : data = 16'b1111101010000110;
            15'b000011111110010 : data = 16'b1111101010001100;
            15'b000011111110011 : data = 16'b1111101010010010;
            15'b000011111110100 : data = 16'b1111101010011000;
            15'b000011111110101 : data = 16'b1111101010011110;
            15'b000011111110110 : data = 16'b1111101010100100;
            15'b000011111110111 : data = 16'b1111101010101010;
            15'b000011111111000 : data = 16'b1111101010101111;
            15'b000011111111001 : data = 16'b1111101010110101;
            15'b000011111111010 : data = 16'b1111101010111011;
            15'b000011111111011 : data = 16'b1111101011000001;
            15'b000011111111100 : data = 16'b1111101011000111;
            15'b000011111111101 : data = 16'b1111101011001101;
            15'b000011111111110 : data = 16'b1111101011010010;
            15'b000011111111111 : data = 16'b1111101011011000;
            15'b000100000000000 : data = 16'b1111101011011110;
            15'b000100000000001 : data = 16'b1111101011100100;
            15'b000100000000010 : data = 16'b1111101011101001;
            15'b000100000000011 : data = 16'b1111101011101111;
            15'b000100000000100 : data = 16'b1111101011110101;
            15'b000100000000101 : data = 16'b1111101011111011;
            15'b000100000000110 : data = 16'b1111101100000000;
            15'b000100000000111 : data = 16'b1111101100000110;
            15'b000100000001000 : data = 16'b1111101100001100;
            15'b000100000001001 : data = 16'b1111101100010001;
            15'b000100000001010 : data = 16'b1111101100010111;
            15'b000100000001011 : data = 16'b1111101100011101;
            15'b000100000001100 : data = 16'b1111101100100010;
            15'b000100000001101 : data = 16'b1111101100101000;
            15'b000100000001110 : data = 16'b1111101100101101;
            15'b000100000001111 : data = 16'b1111101100110011;
            15'b000100000010000 : data = 16'b1111101100111001;
            15'b000100000010001 : data = 16'b1111101100111110;
            15'b000100000010010 : data = 16'b1111101101000100;
            15'b000100000010011 : data = 16'b1111101101001001;
            15'b000100000010100 : data = 16'b1111101101001111;
            15'b000100000010101 : data = 16'b1111101101010100;
            15'b000100000010110 : data = 16'b1111101101011010;
            15'b000100000010111 : data = 16'b1111101101011111;
            15'b000100000011000 : data = 16'b1111101101100101;
            15'b000100000011001 : data = 16'b1111101101101010;
            15'b000100000011010 : data = 16'b1111101101110000;
            15'b000100000011011 : data = 16'b1111101101110101;
            15'b000100000011100 : data = 16'b1111101101111011;
            15'b000100000011101 : data = 16'b1111101110000000;
            15'b000100000011110 : data = 16'b1111101110000101;
            15'b000100000011111 : data = 16'b1111101110001011;
            15'b000100000100000 : data = 16'b1111101110010000;
            15'b000100000100001 : data = 16'b1111101110010110;
            15'b000100000100010 : data = 16'b1111101110011011;
            15'b000100000100011 : data = 16'b1111101110100000;
            15'b000100000100100 : data = 16'b1111101110100110;
            15'b000100000100101 : data = 16'b1111101110101011;
            15'b000100000100110 : data = 16'b1111101110110000;
            15'b000100000100111 : data = 16'b1111101110110101;
            15'b000100000101000 : data = 16'b1111101110111011;
            15'b000100000101001 : data = 16'b1111101111000000;
            15'b000100000101010 : data = 16'b1111101111000101;
            15'b000100000101011 : data = 16'b1111101111001010;
            15'b000100000101100 : data = 16'b1111101111010000;
            15'b000100000101101 : data = 16'b1111101111010101;
            15'b000100000101110 : data = 16'b1111101111011010;
            15'b000100000101111 : data = 16'b1111101111011111;
            15'b000100000110000 : data = 16'b1111101111100100;
            15'b000100000110001 : data = 16'b1111101111101010;
            15'b000100000110010 : data = 16'b1111101111101111;
            15'b000100000110011 : data = 16'b1111101111110100;
            15'b000100000110100 : data = 16'b1111101111111001;
            15'b000100000110101 : data = 16'b1111101111111110;
            15'b000100000110110 : data = 16'b1111110000000011;
            15'b000100000110111 : data = 16'b1111110000001000;
            15'b000100000111000 : data = 16'b1111110000001101;
            15'b000100000111001 : data = 16'b1111110000010011;
            15'b000100000111010 : data = 16'b1111110000011000;
            15'b000100000111011 : data = 16'b1111110000011101;
            15'b000100000111100 : data = 16'b1111110000100010;
            15'b000100000111101 : data = 16'b1111110000100111;
            15'b000100000111110 : data = 16'b1111110000101100;
            15'b000100000111111 : data = 16'b1111110000110001;
            15'b000100001000000 : data = 16'b1111110000110110;
            15'b000100001000001 : data = 16'b1111110000111011;
            15'b000100001000010 : data = 16'b1111110001000000;
            15'b000100001000011 : data = 16'b1111110001000100;
            15'b000100001000100 : data = 16'b1111110001001001;
            15'b000100001000101 : data = 16'b1111110001001110;
            15'b000100001000110 : data = 16'b1111110001010011;
            15'b000100001000111 : data = 16'b1111110001011000;
            15'b000100001001000 : data = 16'b1111110001011101;
            15'b000100001001001 : data = 16'b1111110001100010;
            15'b000100001001010 : data = 16'b1111110001100111;
            15'b000100001001011 : data = 16'b1111110001101100;
            15'b000100001001100 : data = 16'b1111110001110000;
            15'b000100001001101 : data = 16'b1111110001110101;
            15'b000100001001110 : data = 16'b1111110001111010;
            15'b000100001001111 : data = 16'b1111110001111111;
            15'b000100001010000 : data = 16'b1111110010000100;
            15'b000100001010001 : data = 16'b1111110010001000;
            15'b000100001010010 : data = 16'b1111110010001101;
            15'b000100001010011 : data = 16'b1111110010010010;
            15'b000100001010100 : data = 16'b1111110010010110;
            15'b000100001010101 : data = 16'b1111110010011011;
            15'b000100001010110 : data = 16'b1111110010100000;
            15'b000100001010111 : data = 16'b1111110010100101;
            15'b000100001011000 : data = 16'b1111110010101001;
            15'b000100001011001 : data = 16'b1111110010101110;
            15'b000100001011010 : data = 16'b1111110010110011;
            15'b000100001011011 : data = 16'b1111110010110111;
            15'b000100001011100 : data = 16'b1111110010111100;
            15'b000100001011101 : data = 16'b1111110011000000;
            15'b000100001011110 : data = 16'b1111110011000101;
            15'b000100001011111 : data = 16'b1111110011001010;
            15'b000100001100000 : data = 16'b1111110011001110;
            15'b000100001100001 : data = 16'b1111110011010011;
            15'b000100001100010 : data = 16'b1111110011010111;
            15'b000100001100011 : data = 16'b1111110011011100;
            15'b000100001100100 : data = 16'b1111110011100000;
            15'b000100001100101 : data = 16'b1111110011100101;
            15'b000100001100110 : data = 16'b1111110011101001;
            15'b000100001100111 : data = 16'b1111110011101110;
            15'b000100001101000 : data = 16'b1111110011110010;
            15'b000100001101001 : data = 16'b1111110011110111;
            15'b000100001101010 : data = 16'b1111110011111011;
            15'b000100001101011 : data = 16'b1111110100000000;
            15'b000100001101100 : data = 16'b1111110100000100;
            15'b000100001101101 : data = 16'b1111110100001000;
            15'b000100001101110 : data = 16'b1111110100001101;
            15'b000100001101111 : data = 16'b1111110100010001;
            15'b000100001110000 : data = 16'b1111110100010110;
            15'b000100001110001 : data = 16'b1111110100011010;
            15'b000100001110010 : data = 16'b1111110100011110;
            15'b000100001110011 : data = 16'b1111110100100011;
            15'b000100001110100 : data = 16'b1111110100100111;
            15'b000100001110101 : data = 16'b1111110100101011;
            15'b000100001110110 : data = 16'b1111110100110000;
            15'b000100001110111 : data = 16'b1111110100110100;
            15'b000100001111000 : data = 16'b1111110100111000;
            15'b000100001111001 : data = 16'b1111110100111100;
            15'b000100001111010 : data = 16'b1111110101000001;
            15'b000100001111011 : data = 16'b1111110101000101;
            15'b000100001111100 : data = 16'b1111110101001001;
            15'b000100001111101 : data = 16'b1111110101001101;
            15'b000100001111110 : data = 16'b1111110101010010;
            15'b000100001111111 : data = 16'b1111110101010110;
            15'b000100010000000 : data = 16'b1111110101011010;
            15'b000100010000001 : data = 16'b1111110101011110;
            15'b000100010000010 : data = 16'b1111110101100010;
            15'b000100010000011 : data = 16'b1111110101100110;
            15'b000100010000100 : data = 16'b1111110101101010;
            15'b000100010000101 : data = 16'b1111110101101111;
            15'b000100010000110 : data = 16'b1111110101110011;
            15'b000100010000111 : data = 16'b1111110101110111;
            15'b000100010001000 : data = 16'b1111110101111011;
            15'b000100010001001 : data = 16'b1111110101111111;
            15'b000100010001010 : data = 16'b1111110110000011;
            15'b000100010001011 : data = 16'b1111110110000111;
            15'b000100010001100 : data = 16'b1111110110001011;
            15'b000100010001101 : data = 16'b1111110110001111;
            15'b000100010001110 : data = 16'b1111110110010011;
            15'b000100010001111 : data = 16'b1111110110010111;
            15'b000100010010000 : data = 16'b1111110110011011;
            15'b000100010010001 : data = 16'b1111110110011111;
            15'b000100010010010 : data = 16'b1111110110100011;
            15'b000100010010011 : data = 16'b1111110110100111;
            15'b000100010010100 : data = 16'b1111110110101011;
            15'b000100010010101 : data = 16'b1111110110101110;
            15'b000100010010110 : data = 16'b1111110110110010;
            15'b000100010010111 : data = 16'b1111110110110110;
            15'b000100010011000 : data = 16'b1111110110111010;
            15'b000100010011001 : data = 16'b1111110110111110;
            15'b000100010011010 : data = 16'b1111110111000010;
            15'b000100010011011 : data = 16'b1111110111000110;
            15'b000100010011100 : data = 16'b1111110111001001;
            15'b000100010011101 : data = 16'b1111110111001101;
            15'b000100010011110 : data = 16'b1111110111010001;
            15'b000100010011111 : data = 16'b1111110111010101;
            15'b000100010100000 : data = 16'b1111110111011001;
            15'b000100010100001 : data = 16'b1111110111011100;
            15'b000100010100010 : data = 16'b1111110111100000;
            15'b000100010100011 : data = 16'b1111110111100100;
            15'b000100010100100 : data = 16'b1111110111100111;
            15'b000100010100101 : data = 16'b1111110111101011;
            15'b000100010100110 : data = 16'b1111110111101111;
            15'b000100010100111 : data = 16'b1111110111110011;
            15'b000100010101000 : data = 16'b1111110111110110;
            15'b000100010101001 : data = 16'b1111110111111010;
            15'b000100010101010 : data = 16'b1111110111111101;
            15'b000100010101011 : data = 16'b1111111000000001;
            15'b000100010101100 : data = 16'b1111111000000101;
            15'b000100010101101 : data = 16'b1111111000001000;
            15'b000100010101110 : data = 16'b1111111000001100;
            15'b000100010101111 : data = 16'b1111111000001111;
            15'b000100010110000 : data = 16'b1111111000010011;
            15'b000100010110001 : data = 16'b1111111000010111;
            15'b000100010110010 : data = 16'b1111111000011010;
            15'b000100010110011 : data = 16'b1111111000011110;
            15'b000100010110100 : data = 16'b1111111000100001;
            15'b000100010110101 : data = 16'b1111111000100101;
            15'b000100010110110 : data = 16'b1111111000101000;
            15'b000100010110111 : data = 16'b1111111000101100;
            15'b000100010111000 : data = 16'b1111111000101111;
            15'b000100010111001 : data = 16'b1111111000110010;
            15'b000100010111010 : data = 16'b1111111000110110;
            15'b000100010111011 : data = 16'b1111111000111001;
            15'b000100010111100 : data = 16'b1111111000111101;
            15'b000100010111101 : data = 16'b1111111001000000;
            15'b000100010111110 : data = 16'b1111111001000100;
            15'b000100010111111 : data = 16'b1111111001000111;
            15'b000100011000000 : data = 16'b1111111001001010;
            15'b000100011000001 : data = 16'b1111111001001110;
            15'b000100011000010 : data = 16'b1111111001010001;
            15'b000100011000011 : data = 16'b1111111001010100;
            15'b000100011000100 : data = 16'b1111111001011000;
            15'b000100011000101 : data = 16'b1111111001011011;
            15'b000100011000110 : data = 16'b1111111001011110;
            15'b000100011000111 : data = 16'b1111111001100001;
            15'b000100011001000 : data = 16'b1111111001100101;
            15'b000100011001001 : data = 16'b1111111001101000;
            15'b000100011001010 : data = 16'b1111111001101011;
            15'b000100011001011 : data = 16'b1111111001101110;
            15'b000100011001100 : data = 16'b1111111001110001;
            15'b000100011001101 : data = 16'b1111111001110101;
            15'b000100011001110 : data = 16'b1111111001111000;
            15'b000100011001111 : data = 16'b1111111001111011;
            15'b000100011010000 : data = 16'b1111111001111110;
            15'b000100011010001 : data = 16'b1111111010000001;
            15'b000100011010010 : data = 16'b1111111010000100;
            15'b000100011010011 : data = 16'b1111111010001000;
            15'b000100011010100 : data = 16'b1111111010001011;
            15'b000100011010101 : data = 16'b1111111010001110;
            15'b000100011010110 : data = 16'b1111111010010001;
            15'b000100011010111 : data = 16'b1111111010010100;
            15'b000100011011000 : data = 16'b1111111010010111;
            15'b000100011011001 : data = 16'b1111111010011010;
            15'b000100011011010 : data = 16'b1111111010011101;
            15'b000100011011011 : data = 16'b1111111010100000;
            15'b000100011011100 : data = 16'b1111111010100011;
            15'b000100011011101 : data = 16'b1111111010100110;
            15'b000100011011110 : data = 16'b1111111010101001;
            15'b000100011011111 : data = 16'b1111111010101100;
            15'b000100011100000 : data = 16'b1111111010101111;
            15'b000100011100001 : data = 16'b1111111010110010;
            15'b000100011100010 : data = 16'b1111111010110101;
            15'b000100011100011 : data = 16'b1111111010111000;
            15'b000100011100100 : data = 16'b1111111010111010;
            15'b000100011100101 : data = 16'b1111111010111101;
            15'b000100011100110 : data = 16'b1111111011000000;
            15'b000100011100111 : data = 16'b1111111011000011;
            15'b000100011101000 : data = 16'b1111111011000110;
            15'b000100011101001 : data = 16'b1111111011001001;
            15'b000100011101010 : data = 16'b1111111011001100;
            15'b000100011101011 : data = 16'b1111111011001110;
            15'b000100011101100 : data = 16'b1111111011010001;
            15'b000100011101101 : data = 16'b1111111011010100;
            15'b000100011101110 : data = 16'b1111111011010111;
            15'b000100011101111 : data = 16'b1111111011011001;
            15'b000100011110000 : data = 16'b1111111011011100;
            15'b000100011110001 : data = 16'b1111111011011111;
            15'b000100011110010 : data = 16'b1111111011100010;
            15'b000100011110011 : data = 16'b1111111011100100;
            15'b000100011110100 : data = 16'b1111111011100111;
            15'b000100011110101 : data = 16'b1111111011101010;
            15'b000100011110110 : data = 16'b1111111011101100;
            15'b000100011110111 : data = 16'b1111111011101111;
            15'b000100011111000 : data = 16'b1111111011110010;
            15'b000100011111001 : data = 16'b1111111011110100;
            15'b000100011111010 : data = 16'b1111111011110111;
            15'b000100011111011 : data = 16'b1111111011111010;
            15'b000100011111100 : data = 16'b1111111011111100;
            15'b000100011111101 : data = 16'b1111111011111111;
            15'b000100011111110 : data = 16'b1111111100000001;
            15'b000100011111111 : data = 16'b1111111100000100;
            15'b000100100000000 : data = 16'b1111111100000110;
            15'b000100100000001 : data = 16'b1111111100001001;
            15'b000100100000010 : data = 16'b1111111100001011;
            15'b000100100000011 : data = 16'b1111111100001110;
            15'b000100100000100 : data = 16'b1111111100010000;
            15'b000100100000101 : data = 16'b1111111100010011;
            15'b000100100000110 : data = 16'b1111111100010101;
            15'b000100100000111 : data = 16'b1111111100011000;
            15'b000100100001000 : data = 16'b1111111100011010;
            15'b000100100001001 : data = 16'b1111111100011101;
            15'b000100100001010 : data = 16'b1111111100011111;
            15'b000100100001011 : data = 16'b1111111100100001;
            15'b000100100001100 : data = 16'b1111111100100100;
            15'b000100100001101 : data = 16'b1111111100100110;
            15'b000100100001110 : data = 16'b1111111100101000;
            15'b000100100001111 : data = 16'b1111111100101011;
            15'b000100100010000 : data = 16'b1111111100101101;
            15'b000100100010001 : data = 16'b1111111100101111;
            15'b000100100010010 : data = 16'b1111111100110010;
            15'b000100100010011 : data = 16'b1111111100110100;
            15'b000100100010100 : data = 16'b1111111100110110;
            15'b000100100010101 : data = 16'b1111111100111001;
            15'b000100100010110 : data = 16'b1111111100111011;
            15'b000100100010111 : data = 16'b1111111100111101;
            15'b000100100011000 : data = 16'b1111111100111111;
            15'b000100100011001 : data = 16'b1111111101000010;
            15'b000100100011010 : data = 16'b1111111101000100;
            15'b000100100011011 : data = 16'b1111111101000110;
            15'b000100100011100 : data = 16'b1111111101001000;
            15'b000100100011101 : data = 16'b1111111101001010;
            15'b000100100011110 : data = 16'b1111111101001100;
            15'b000100100011111 : data = 16'b1111111101001111;
            15'b000100100100000 : data = 16'b1111111101010001;
            15'b000100100100001 : data = 16'b1111111101010011;
            15'b000100100100010 : data = 16'b1111111101010101;
            15'b000100100100011 : data = 16'b1111111101010111;
            15'b000100100100100 : data = 16'b1111111101011001;
            15'b000100100100101 : data = 16'b1111111101011011;
            15'b000100100100110 : data = 16'b1111111101011101;
            15'b000100100100111 : data = 16'b1111111101011111;
            15'b000100100101000 : data = 16'b1111111101100001;
            15'b000100100101001 : data = 16'b1111111101100011;
            15'b000100100101010 : data = 16'b1111111101100101;
            15'b000100100101011 : data = 16'b1111111101100111;
            15'b000100100101100 : data = 16'b1111111101101001;
            15'b000100100101101 : data = 16'b1111111101101011;
            15'b000100100101110 : data = 16'b1111111101101101;
            15'b000100100101111 : data = 16'b1111111101101111;
            15'b000100100110000 : data = 16'b1111111101110001;
            15'b000100100110001 : data = 16'b1111111101110011;
            15'b000100100110010 : data = 16'b1111111101110101;
            15'b000100100110011 : data = 16'b1111111101110111;
            15'b000100100110100 : data = 16'b1111111101111000;
            15'b000100100110101 : data = 16'b1111111101111010;
            15'b000100100110110 : data = 16'b1111111101111100;
            15'b000100100110111 : data = 16'b1111111101111110;
            15'b000100100111000 : data = 16'b1111111110000000;
            15'b000100100111001 : data = 16'b1111111110000010;
            15'b000100100111010 : data = 16'b1111111110000011;
            15'b000100100111011 : data = 16'b1111111110000101;
            15'b000100100111100 : data = 16'b1111111110000111;
            15'b000100100111101 : data = 16'b1111111110001001;
            15'b000100100111110 : data = 16'b1111111110001010;
            15'b000100100111111 : data = 16'b1111111110001100;
            15'b000100101000000 : data = 16'b1111111110001110;
            15'b000100101000001 : data = 16'b1111111110010000;
            15'b000100101000010 : data = 16'b1111111110010001;
            15'b000100101000011 : data = 16'b1111111110010011;
            15'b000100101000100 : data = 16'b1111111110010101;
            15'b000100101000101 : data = 16'b1111111110010110;
            15'b000100101000110 : data = 16'b1111111110011000;
            15'b000100101000111 : data = 16'b1111111110011001;
            15'b000100101001000 : data = 16'b1111111110011011;
            15'b000100101001001 : data = 16'b1111111110011101;
            15'b000100101001010 : data = 16'b1111111110011110;
            15'b000100101001011 : data = 16'b1111111110100000;
            15'b000100101001100 : data = 16'b1111111110100001;
            15'b000100101001101 : data = 16'b1111111110100011;
            15'b000100101001110 : data = 16'b1111111110100100;
            15'b000100101001111 : data = 16'b1111111110100110;
            15'b000100101010000 : data = 16'b1111111110101000;
            15'b000100101010001 : data = 16'b1111111110101001;
            15'b000100101010010 : data = 16'b1111111110101010;
            15'b000100101010011 : data = 16'b1111111110101100;
            15'b000100101010100 : data = 16'b1111111110101101;
            15'b000100101010101 : data = 16'b1111111110101111;
            15'b000100101010110 : data = 16'b1111111110110000;
            15'b000100101010111 : data = 16'b1111111110110010;
            15'b000100101011000 : data = 16'b1111111110110011;
            15'b000100101011001 : data = 16'b1111111110110100;
            15'b000100101011010 : data = 16'b1111111110110110;
            15'b000100101011011 : data = 16'b1111111110110111;
            15'b000100101011100 : data = 16'b1111111110111001;
            15'b000100101011101 : data = 16'b1111111110111010;
            15'b000100101011110 : data = 16'b1111111110111011;
            15'b000100101011111 : data = 16'b1111111110111101;
            15'b000100101100000 : data = 16'b1111111110111110;
            15'b000100101100001 : data = 16'b1111111110111111;
            15'b000100101100010 : data = 16'b1111111111000000;
            15'b000100101100011 : data = 16'b1111111111000010;
            15'b000100101100100 : data = 16'b1111111111000011;
            15'b000100101100101 : data = 16'b1111111111000100;
            15'b000100101100110 : data = 16'b1111111111000101;
            15'b000100101100111 : data = 16'b1111111111000111;
            15'b000100101101000 : data = 16'b1111111111001000;
            15'b000100101101001 : data = 16'b1111111111001001;
            15'b000100101101010 : data = 16'b1111111111001010;
            15'b000100101101011 : data = 16'b1111111111001011;
            15'b000100101101100 : data = 16'b1111111111001100;
            15'b000100101101101 : data = 16'b1111111111001110;
            15'b000100101101110 : data = 16'b1111111111001111;
            15'b000100101101111 : data = 16'b1111111111010000;
            15'b000100101110000 : data = 16'b1111111111010001;
            15'b000100101110001 : data = 16'b1111111111010010;
            15'b000100101110010 : data = 16'b1111111111010011;
            15'b000100101110011 : data = 16'b1111111111010100;
            15'b000100101110100 : data = 16'b1111111111010101;
            15'b000100101110101 : data = 16'b1111111111010110;
            15'b000100101110110 : data = 16'b1111111111010111;
            15'b000100101110111 : data = 16'b1111111111011000;
            15'b000100101111000 : data = 16'b1111111111011001;
            15'b000100101111001 : data = 16'b1111111111011010;
            15'b000100101111010 : data = 16'b1111111111011011;
            15'b000100101111011 : data = 16'b1111111111011100;
            15'b000100101111100 : data = 16'b1111111111011101;
            15'b000100101111101 : data = 16'b1111111111011110;
            15'b000100101111110 : data = 16'b1111111111011111;
            15'b000100101111111 : data = 16'b1111111111100000;
            15'b000100110000000 : data = 16'b1111111111100001;
            15'b000100110000001 : data = 16'b1111111111100001;
            15'b000100110000010 : data = 16'b1111111111100010;
            15'b000100110000011 : data = 16'b1111111111100011;
            15'b000100110000100 : data = 16'b1111111111100100;
            15'b000100110000101 : data = 16'b1111111111100101;
            15'b000100110000110 : data = 16'b1111111111100110;
            15'b000100110000111 : data = 16'b1111111111100110;
            15'b000100110001000 : data = 16'b1111111111100111;
            15'b000100110001001 : data = 16'b1111111111101000;
            15'b000100110001010 : data = 16'b1111111111101001;
            15'b000100110001011 : data = 16'b1111111111101001;
            15'b000100110001100 : data = 16'b1111111111101010;
            15'b000100110001101 : data = 16'b1111111111101011;
            15'b000100110001110 : data = 16'b1111111111101100;
            15'b000100110001111 : data = 16'b1111111111101100;
            15'b000100110010000 : data = 16'b1111111111101101;
            15'b000100110010001 : data = 16'b1111111111101110;
            15'b000100110010010 : data = 16'b1111111111101110;
            15'b000100110010011 : data = 16'b1111111111101111;
            15'b000100110010100 : data = 16'b1111111111110000;
            15'b000100110010101 : data = 16'b1111111111110000;
            15'b000100110010110 : data = 16'b1111111111110001;
            15'b000100110010111 : data = 16'b1111111111110001;
            15'b000100110011000 : data = 16'b1111111111110010;
            15'b000100110011001 : data = 16'b1111111111110011;
            15'b000100110011010 : data = 16'b1111111111110011;
            15'b000100110011011 : data = 16'b1111111111110100;
            15'b000100110011100 : data = 16'b1111111111110100;
            15'b000100110011101 : data = 16'b1111111111110101;
            15'b000100110011110 : data = 16'b1111111111110101;
            15'b000100110011111 : data = 16'b1111111111110110;
            15'b000100110100000 : data = 16'b1111111111110110;
            15'b000100110100001 : data = 16'b1111111111110111;
            15'b000100110100010 : data = 16'b1111111111110111;
            15'b000100110100011 : data = 16'b1111111111110111;
            15'b000100110100100 : data = 16'b1111111111111000;
            15'b000100110100101 : data = 16'b1111111111111000;
            15'b000100110100110 : data = 16'b1111111111111001;
            15'b000100110100111 : data = 16'b1111111111111001;
            15'b000100110101000 : data = 16'b1111111111111001;
            15'b000100110101001 : data = 16'b1111111111111010;
            15'b000100110101010 : data = 16'b1111111111111010;
            15'b000100110101011 : data = 16'b1111111111111010;
            15'b000100110101100 : data = 16'b1111111111111011;
            15'b000100110101101 : data = 16'b1111111111111011;
            15'b000100110101110 : data = 16'b1111111111111011;
            15'b000100110101111 : data = 16'b1111111111111100;
            15'b000100110110000 : data = 16'b1111111111111100;
            15'b000100110110001 : data = 16'b1111111111111100;
            15'b000100110110010 : data = 16'b1111111111111100;
            15'b000100110110011 : data = 16'b1111111111111101;
            15'b000100110110100 : data = 16'b1111111111111101;
            15'b000100110110101 : data = 16'b1111111111111101;
            15'b000100110110110 : data = 16'b1111111111111101;
            15'b000100110110111 : data = 16'b1111111111111101;
            15'b000100110111000 : data = 16'b1111111111111110;
            15'b000100110111001 : data = 16'b1111111111111110;
            15'b000100110111010 : data = 16'b1111111111111110;
            15'b000100110111011 : data = 16'b1111111111111110;
            15'b000100110111100 : data = 16'b1111111111111110;
            15'b000100110111101 : data = 16'b1111111111111110;
            15'b000100110111110 : data = 16'b1111111111111110;
            15'b000100110111111 : data = 16'b1111111111111110;
            15'b000100111000000 : data = 16'b1111111111111110;
            15'b000100111000001 : data = 16'b1111111111111110;
            15'b000100111000010 : data = 16'b1111111111111110;
            15'b000100111000011 : data = 16'b1111111111111110;
            15'b000100111000100 : data = 16'b1111111111111111;
            15'b000100111000101 : data = 16'b1111111111111110;
            15'b000100111000110 : data = 16'b1111111111111110;
            15'b000100111000111 : data = 16'b1111111111111110;
            15'b000100111001000 : data = 16'b1111111111111110;
            15'b000100111001001 : data = 16'b1111111111111110;
            15'b000100111001010 : data = 16'b1111111111111110;
            15'b000100111001011 : data = 16'b1111111111111110;
            15'b000100111001100 : data = 16'b1111111111111110;
            15'b000100111001101 : data = 16'b1111111111111110;
            15'b000100111001110 : data = 16'b1111111111111110;
            15'b000100111001111 : data = 16'b1111111111111110;
            15'b000100111010000 : data = 16'b1111111111111110;
            15'b000100111010001 : data = 16'b1111111111111101;
            15'b000100111010010 : data = 16'b1111111111111101;
            15'b000100111010011 : data = 16'b1111111111111101;
            15'b000100111010100 : data = 16'b1111111111111101;
            15'b000100111010101 : data = 16'b1111111111111101;
            15'b000100111010110 : data = 16'b1111111111111100;
            15'b000100111010111 : data = 16'b1111111111111100;
            15'b000100111011000 : data = 16'b1111111111111100;
            15'b000100111011001 : data = 16'b1111111111111100;
            15'b000100111011010 : data = 16'b1111111111111011;
            15'b000100111011011 : data = 16'b1111111111111011;
            15'b000100111011100 : data = 16'b1111111111111011;
            15'b000100111011101 : data = 16'b1111111111111010;
            15'b000100111011110 : data = 16'b1111111111111010;
            15'b000100111011111 : data = 16'b1111111111111010;
            15'b000100111100000 : data = 16'b1111111111111001;
            15'b000100111100001 : data = 16'b1111111111111001;
            15'b000100111100010 : data = 16'b1111111111111001;
            15'b000100111100011 : data = 16'b1111111111111000;
            15'b000100111100100 : data = 16'b1111111111111000;
            15'b000100111100101 : data = 16'b1111111111110111;
            15'b000100111100110 : data = 16'b1111111111110111;
            15'b000100111100111 : data = 16'b1111111111110111;
            15'b000100111101000 : data = 16'b1111111111110110;
            15'b000100111101001 : data = 16'b1111111111110110;
            15'b000100111101010 : data = 16'b1111111111110101;
            15'b000100111101011 : data = 16'b1111111111110101;
            15'b000100111101100 : data = 16'b1111111111110100;
            15'b000100111101101 : data = 16'b1111111111110100;
            15'b000100111101110 : data = 16'b1111111111110011;
            15'b000100111101111 : data = 16'b1111111111110011;
            15'b000100111110000 : data = 16'b1111111111110010;
            15'b000100111110001 : data = 16'b1111111111110001;
            15'b000100111110010 : data = 16'b1111111111110001;
            15'b000100111110011 : data = 16'b1111111111110000;
            15'b000100111110100 : data = 16'b1111111111110000;
            15'b000100111110101 : data = 16'b1111111111101111;
            15'b000100111110110 : data = 16'b1111111111101110;
            15'b000100111110111 : data = 16'b1111111111101110;
            15'b000100111111000 : data = 16'b1111111111101101;
            15'b000100111111001 : data = 16'b1111111111101100;
            15'b000100111111010 : data = 16'b1111111111101100;
            15'b000100111111011 : data = 16'b1111111111101011;
            15'b000100111111100 : data = 16'b1111111111101010;
            15'b000100111111101 : data = 16'b1111111111101001;
            15'b000100111111110 : data = 16'b1111111111101001;
            15'b000100111111111 : data = 16'b1111111111101000;
            15'b000101000000000 : data = 16'b1111111111100111;
            15'b000101000000001 : data = 16'b1111111111100110;
            15'b000101000000010 : data = 16'b1111111111100110;
            15'b000101000000011 : data = 16'b1111111111100101;
            15'b000101000000100 : data = 16'b1111111111100100;
            15'b000101000000101 : data = 16'b1111111111100011;
            15'b000101000000110 : data = 16'b1111111111100010;
            15'b000101000000111 : data = 16'b1111111111100001;
            15'b000101000001000 : data = 16'b1111111111100001;
            15'b000101000001001 : data = 16'b1111111111100000;
            15'b000101000001010 : data = 16'b1111111111011111;
            15'b000101000001011 : data = 16'b1111111111011110;
            15'b000101000001100 : data = 16'b1111111111011101;
            15'b000101000001101 : data = 16'b1111111111011100;
            15'b000101000001110 : data = 16'b1111111111011011;
            15'b000101000001111 : data = 16'b1111111111011010;
            15'b000101000010000 : data = 16'b1111111111011001;
            15'b000101000010001 : data = 16'b1111111111011000;
            15'b000101000010010 : data = 16'b1111111111010111;
            15'b000101000010011 : data = 16'b1111111111010110;
            15'b000101000010100 : data = 16'b1111111111010101;
            15'b000101000010101 : data = 16'b1111111111010100;
            15'b000101000010110 : data = 16'b1111111111010011;
            15'b000101000010111 : data = 16'b1111111111010010;
            15'b000101000011000 : data = 16'b1111111111010001;
            15'b000101000011001 : data = 16'b1111111111010000;
            15'b000101000011010 : data = 16'b1111111111001111;
            15'b000101000011011 : data = 16'b1111111111001110;
            15'b000101000011100 : data = 16'b1111111111001100;
            15'b000101000011101 : data = 16'b1111111111001011;
            15'b000101000011110 : data = 16'b1111111111001010;
            15'b000101000011111 : data = 16'b1111111111001001;
            15'b000101000100000 : data = 16'b1111111111001000;
            15'b000101000100001 : data = 16'b1111111111000111;
            15'b000101000100010 : data = 16'b1111111111000101;
            15'b000101000100011 : data = 16'b1111111111000100;
            15'b000101000100100 : data = 16'b1111111111000011;
            15'b000101000100101 : data = 16'b1111111111000010;
            15'b000101000100110 : data = 16'b1111111111000000;
            15'b000101000100111 : data = 16'b1111111110111111;
            15'b000101000101000 : data = 16'b1111111110111110;
            15'b000101000101001 : data = 16'b1111111110111101;
            15'b000101000101010 : data = 16'b1111111110111011;
            15'b000101000101011 : data = 16'b1111111110111010;
            15'b000101000101100 : data = 16'b1111111110111001;
            15'b000101000101101 : data = 16'b1111111110110111;
            15'b000101000101110 : data = 16'b1111111110110110;
            15'b000101000101111 : data = 16'b1111111110110100;
            15'b000101000110000 : data = 16'b1111111110110011;
            15'b000101000110001 : data = 16'b1111111110110010;
            15'b000101000110010 : data = 16'b1111111110110000;
            15'b000101000110011 : data = 16'b1111111110101111;
            15'b000101000110100 : data = 16'b1111111110101101;
            15'b000101000110101 : data = 16'b1111111110101100;
            15'b000101000110110 : data = 16'b1111111110101010;
            15'b000101000110111 : data = 16'b1111111110101001;
            15'b000101000111000 : data = 16'b1111111110101000;
            15'b000101000111001 : data = 16'b1111111110100110;
            15'b000101000111010 : data = 16'b1111111110100100;
            15'b000101000111011 : data = 16'b1111111110100011;
            15'b000101000111100 : data = 16'b1111111110100001;
            15'b000101000111101 : data = 16'b1111111110100000;
            15'b000101000111110 : data = 16'b1111111110011110;
            15'b000101000111111 : data = 16'b1111111110011101;
            15'b000101001000000 : data = 16'b1111111110011011;
            15'b000101001000001 : data = 16'b1111111110011001;
            15'b000101001000010 : data = 16'b1111111110011000;
            15'b000101001000011 : data = 16'b1111111110010110;
            15'b000101001000100 : data = 16'b1111111110010101;
            15'b000101001000101 : data = 16'b1111111110010011;
            15'b000101001000110 : data = 16'b1111111110010001;
            15'b000101001000111 : data = 16'b1111111110010000;
            15'b000101001001000 : data = 16'b1111111110001110;
            15'b000101001001001 : data = 16'b1111111110001100;
            15'b000101001001010 : data = 16'b1111111110001010;
            15'b000101001001011 : data = 16'b1111111110001001;
            15'b000101001001100 : data = 16'b1111111110000111;
            15'b000101001001101 : data = 16'b1111111110000101;
            15'b000101001001110 : data = 16'b1111111110000011;
            15'b000101001001111 : data = 16'b1111111110000010;
            15'b000101001010000 : data = 16'b1111111110000000;
            15'b000101001010001 : data = 16'b1111111101111110;
            15'b000101001010010 : data = 16'b1111111101111100;
            15'b000101001010011 : data = 16'b1111111101111010;
            15'b000101001010100 : data = 16'b1111111101111000;
            15'b000101001010101 : data = 16'b1111111101110111;
            15'b000101001010110 : data = 16'b1111111101110101;
            15'b000101001010111 : data = 16'b1111111101110011;
            15'b000101001011000 : data = 16'b1111111101110001;
            15'b000101001011001 : data = 16'b1111111101101111;
            15'b000101001011010 : data = 16'b1111111101101101;
            15'b000101001011011 : data = 16'b1111111101101011;
            15'b000101001011100 : data = 16'b1111111101101001;
            15'b000101001011101 : data = 16'b1111111101100111;
            15'b000101001011110 : data = 16'b1111111101100101;
            15'b000101001011111 : data = 16'b1111111101100011;
            15'b000101001100000 : data = 16'b1111111101100001;
            15'b000101001100001 : data = 16'b1111111101011111;
            15'b000101001100010 : data = 16'b1111111101011101;
            15'b000101001100011 : data = 16'b1111111101011011;
            15'b000101001100100 : data = 16'b1111111101011001;
            15'b000101001100101 : data = 16'b1111111101010111;
            15'b000101001100110 : data = 16'b1111111101010101;
            15'b000101001100111 : data = 16'b1111111101010011;
            15'b000101001101000 : data = 16'b1111111101010001;
            15'b000101001101001 : data = 16'b1111111101001111;
            15'b000101001101010 : data = 16'b1111111101001100;
            15'b000101001101011 : data = 16'b1111111101001010;
            15'b000101001101100 : data = 16'b1111111101001000;
            15'b000101001101101 : data = 16'b1111111101000110;
            15'b000101001101110 : data = 16'b1111111101000100;
            15'b000101001101111 : data = 16'b1111111101000010;
            15'b000101001110000 : data = 16'b1111111100111111;
            15'b000101001110001 : data = 16'b1111111100111101;
            15'b000101001110010 : data = 16'b1111111100111011;
            15'b000101001110011 : data = 16'b1111111100111001;
            15'b000101001110100 : data = 16'b1111111100110110;
            15'b000101001110101 : data = 16'b1111111100110100;
            15'b000101001110110 : data = 16'b1111111100110010;
            15'b000101001110111 : data = 16'b1111111100101111;
            15'b000101001111000 : data = 16'b1111111100101101;
            15'b000101001111001 : data = 16'b1111111100101011;
            15'b000101001111010 : data = 16'b1111111100101000;
            15'b000101001111011 : data = 16'b1111111100100110;
            15'b000101001111100 : data = 16'b1111111100100100;
            15'b000101001111101 : data = 16'b1111111100100001;
            15'b000101001111110 : data = 16'b1111111100011111;
            15'b000101001111111 : data = 16'b1111111100011101;
            15'b000101010000000 : data = 16'b1111111100011010;
            15'b000101010000001 : data = 16'b1111111100011000;
            15'b000101010000010 : data = 16'b1111111100010101;
            15'b000101010000011 : data = 16'b1111111100010011;
            15'b000101010000100 : data = 16'b1111111100010000;
            15'b000101010000101 : data = 16'b1111111100001110;
            15'b000101010000110 : data = 16'b1111111100001011;
            15'b000101010000111 : data = 16'b1111111100001001;
            15'b000101010001000 : data = 16'b1111111100000110;
            15'b000101010001001 : data = 16'b1111111100000100;
            15'b000101010001010 : data = 16'b1111111100000001;
            15'b000101010001011 : data = 16'b1111111011111111;
            15'b000101010001100 : data = 16'b1111111011111100;
            15'b000101010001101 : data = 16'b1111111011111010;
            15'b000101010001110 : data = 16'b1111111011110111;
            15'b000101010001111 : data = 16'b1111111011110100;
            15'b000101010010000 : data = 16'b1111111011110010;
            15'b000101010010001 : data = 16'b1111111011101111;
            15'b000101010010010 : data = 16'b1111111011101100;
            15'b000101010010011 : data = 16'b1111111011101010;
            15'b000101010010100 : data = 16'b1111111011100111;
            15'b000101010010101 : data = 16'b1111111011100100;
            15'b000101010010110 : data = 16'b1111111011100010;
            15'b000101010010111 : data = 16'b1111111011011111;
            15'b000101010011000 : data = 16'b1111111011011100;
            15'b000101010011001 : data = 16'b1111111011011001;
            15'b000101010011010 : data = 16'b1111111011010111;
            15'b000101010011011 : data = 16'b1111111011010100;
            15'b000101010011100 : data = 16'b1111111011010001;
            15'b000101010011101 : data = 16'b1111111011001110;
            15'b000101010011110 : data = 16'b1111111011001100;
            15'b000101010011111 : data = 16'b1111111011001001;
            15'b000101010100000 : data = 16'b1111111011000110;
            15'b000101010100001 : data = 16'b1111111011000011;
            15'b000101010100010 : data = 16'b1111111011000000;
            15'b000101010100011 : data = 16'b1111111010111101;
            15'b000101010100100 : data = 16'b1111111010111010;
            15'b000101010100101 : data = 16'b1111111010111000;
            15'b000101010100110 : data = 16'b1111111010110101;
            15'b000101010100111 : data = 16'b1111111010110010;
            15'b000101010101000 : data = 16'b1111111010101111;
            15'b000101010101001 : data = 16'b1111111010101100;
            15'b000101010101010 : data = 16'b1111111010101001;
            15'b000101010101011 : data = 16'b1111111010100110;
            15'b000101010101100 : data = 16'b1111111010100011;
            15'b000101010101101 : data = 16'b1111111010100000;
            15'b000101010101110 : data = 16'b1111111010011101;
            15'b000101010101111 : data = 16'b1111111010011010;
            15'b000101010110000 : data = 16'b1111111010010111;
            15'b000101010110001 : data = 16'b1111111010010100;
            15'b000101010110010 : data = 16'b1111111010010001;
            15'b000101010110011 : data = 16'b1111111010001110;
            15'b000101010110100 : data = 16'b1111111010001011;
            15'b000101010110101 : data = 16'b1111111010001000;
            15'b000101010110110 : data = 16'b1111111010000100;
            15'b000101010110111 : data = 16'b1111111010000001;
            15'b000101010111000 : data = 16'b1111111001111110;
            15'b000101010111001 : data = 16'b1111111001111011;
            15'b000101010111010 : data = 16'b1111111001111000;
            15'b000101010111011 : data = 16'b1111111001110101;
            15'b000101010111100 : data = 16'b1111111001110001;
            15'b000101010111101 : data = 16'b1111111001101110;
            15'b000101010111110 : data = 16'b1111111001101011;
            15'b000101010111111 : data = 16'b1111111001101000;
            15'b000101011000000 : data = 16'b1111111001100101;
            15'b000101011000001 : data = 16'b1111111001100001;
            15'b000101011000010 : data = 16'b1111111001011110;
            15'b000101011000011 : data = 16'b1111111001011011;
            15'b000101011000100 : data = 16'b1111111001011000;
            15'b000101011000101 : data = 16'b1111111001010100;
            15'b000101011000110 : data = 16'b1111111001010001;
            15'b000101011000111 : data = 16'b1111111001001110;
            15'b000101011001000 : data = 16'b1111111001001010;
            15'b000101011001001 : data = 16'b1111111001000111;
            15'b000101011001010 : data = 16'b1111111001000100;
            15'b000101011001011 : data = 16'b1111111001000000;
            15'b000101011001100 : data = 16'b1111111000111101;
            15'b000101011001101 : data = 16'b1111111000111001;
            15'b000101011001110 : data = 16'b1111111000110110;
            15'b000101011001111 : data = 16'b1111111000110010;
            15'b000101011010000 : data = 16'b1111111000101111;
            15'b000101011010001 : data = 16'b1111111000101100;
            15'b000101011010010 : data = 16'b1111111000101000;
            15'b000101011010011 : data = 16'b1111111000100101;
            15'b000101011010100 : data = 16'b1111111000100001;
            15'b000101011010101 : data = 16'b1111111000011110;
            15'b000101011010110 : data = 16'b1111111000011010;
            15'b000101011010111 : data = 16'b1111111000010111;
            15'b000101011011000 : data = 16'b1111111000010011;
            15'b000101011011001 : data = 16'b1111111000001111;
            15'b000101011011010 : data = 16'b1111111000001100;
            15'b000101011011011 : data = 16'b1111111000001000;
            15'b000101011011100 : data = 16'b1111111000000101;
            15'b000101011011101 : data = 16'b1111111000000001;
            15'b000101011011110 : data = 16'b1111110111111101;
            15'b000101011011111 : data = 16'b1111110111111010;
            15'b000101011100000 : data = 16'b1111110111110110;
            15'b000101011100001 : data = 16'b1111110111110011;
            15'b000101011100010 : data = 16'b1111110111101111;
            15'b000101011100011 : data = 16'b1111110111101011;
            15'b000101011100100 : data = 16'b1111110111100111;
            15'b000101011100101 : data = 16'b1111110111100100;
            15'b000101011100110 : data = 16'b1111110111100000;
            15'b000101011100111 : data = 16'b1111110111011100;
            15'b000101011101000 : data = 16'b1111110111011001;
            15'b000101011101001 : data = 16'b1111110111010101;
            15'b000101011101010 : data = 16'b1111110111010001;
            15'b000101011101011 : data = 16'b1111110111001101;
            15'b000101011101100 : data = 16'b1111110111001001;
            15'b000101011101101 : data = 16'b1111110111000110;
            15'b000101011101110 : data = 16'b1111110111000010;
            15'b000101011101111 : data = 16'b1111110110111110;
            15'b000101011110000 : data = 16'b1111110110111010;
            15'b000101011110001 : data = 16'b1111110110110110;
            15'b000101011110010 : data = 16'b1111110110110010;
            15'b000101011110011 : data = 16'b1111110110101110;
            15'b000101011110100 : data = 16'b1111110110101011;
            15'b000101011110101 : data = 16'b1111110110100111;
            15'b000101011110110 : data = 16'b1111110110100011;
            15'b000101011110111 : data = 16'b1111110110011111;
            15'b000101011111000 : data = 16'b1111110110011011;
            15'b000101011111001 : data = 16'b1111110110010111;
            15'b000101011111010 : data = 16'b1111110110010011;
            15'b000101011111011 : data = 16'b1111110110001111;
            15'b000101011111100 : data = 16'b1111110110001011;
            15'b000101011111101 : data = 16'b1111110110000111;
            15'b000101011111110 : data = 16'b1111110110000011;
            15'b000101011111111 : data = 16'b1111110101111111;
            15'b000101100000000 : data = 16'b1111110101111011;
            15'b000101100000001 : data = 16'b1111110101110111;
            15'b000101100000010 : data = 16'b1111110101110011;
            15'b000101100000011 : data = 16'b1111110101101111;
            15'b000101100000100 : data = 16'b1111110101101010;
            15'b000101100000101 : data = 16'b1111110101100110;
            15'b000101100000110 : data = 16'b1111110101100010;
            15'b000101100000111 : data = 16'b1111110101011110;
            15'b000101100001000 : data = 16'b1111110101011010;
            15'b000101100001001 : data = 16'b1111110101010110;
            15'b000101100001010 : data = 16'b1111110101010010;
            15'b000101100001011 : data = 16'b1111110101001101;
            15'b000101100001100 : data = 16'b1111110101001001;
            15'b000101100001101 : data = 16'b1111110101000101;
            15'b000101100001110 : data = 16'b1111110101000001;
            15'b000101100001111 : data = 16'b1111110100111100;
            15'b000101100010000 : data = 16'b1111110100111000;
            15'b000101100010001 : data = 16'b1111110100110100;
            15'b000101100010010 : data = 16'b1111110100110000;
            15'b000101100010011 : data = 16'b1111110100101011;
            15'b000101100010100 : data = 16'b1111110100100111;
            15'b000101100010101 : data = 16'b1111110100100011;
            15'b000101100010110 : data = 16'b1111110100011110;
            15'b000101100010111 : data = 16'b1111110100011010;
            15'b000101100011000 : data = 16'b1111110100010110;
            15'b000101100011001 : data = 16'b1111110100010001;
            15'b000101100011010 : data = 16'b1111110100001101;
            15'b000101100011011 : data = 16'b1111110100001000;
            15'b000101100011100 : data = 16'b1111110100000100;
            15'b000101100011101 : data = 16'b1111110100000000;
            15'b000101100011110 : data = 16'b1111110011111011;
            15'b000101100011111 : data = 16'b1111110011110111;
            15'b000101100100000 : data = 16'b1111110011110010;
            15'b000101100100001 : data = 16'b1111110011101110;
            15'b000101100100010 : data = 16'b1111110011101001;
            15'b000101100100011 : data = 16'b1111110011100101;
            15'b000101100100100 : data = 16'b1111110011100000;
            15'b000101100100101 : data = 16'b1111110011011100;
            15'b000101100100110 : data = 16'b1111110011010111;
            15'b000101100100111 : data = 16'b1111110011010011;
            15'b000101100101000 : data = 16'b1111110011001110;
            15'b000101100101001 : data = 16'b1111110011001010;
            15'b000101100101010 : data = 16'b1111110011000101;
            15'b000101100101011 : data = 16'b1111110011000000;
            15'b000101100101100 : data = 16'b1111110010111100;
            15'b000101100101101 : data = 16'b1111110010110111;
            15'b000101100101110 : data = 16'b1111110010110011;
            15'b000101100101111 : data = 16'b1111110010101110;
            15'b000101100110000 : data = 16'b1111110010101001;
            15'b000101100110001 : data = 16'b1111110010100101;
            15'b000101100110010 : data = 16'b1111110010100000;
            15'b000101100110011 : data = 16'b1111110010011011;
            15'b000101100110100 : data = 16'b1111110010010110;
            15'b000101100110101 : data = 16'b1111110010010010;
            15'b000101100110110 : data = 16'b1111110010001101;
            15'b000101100110111 : data = 16'b1111110010001000;
            15'b000101100111000 : data = 16'b1111110010000100;
            15'b000101100111001 : data = 16'b1111110001111111;
            15'b000101100111010 : data = 16'b1111110001111010;
            15'b000101100111011 : data = 16'b1111110001110101;
            15'b000101100111100 : data = 16'b1111110001110000;
            15'b000101100111101 : data = 16'b1111110001101100;
            15'b000101100111110 : data = 16'b1111110001100111;
            15'b000101100111111 : data = 16'b1111110001100010;
            15'b000101101000000 : data = 16'b1111110001011101;
            15'b000101101000001 : data = 16'b1111110001011000;
            15'b000101101000010 : data = 16'b1111110001010011;
            15'b000101101000011 : data = 16'b1111110001001110;
            15'b000101101000100 : data = 16'b1111110001001001;
            15'b000101101000101 : data = 16'b1111110001000100;
            15'b000101101000110 : data = 16'b1111110001000000;
            15'b000101101000111 : data = 16'b1111110000111011;
            15'b000101101001000 : data = 16'b1111110000110110;
            15'b000101101001001 : data = 16'b1111110000110001;
            15'b000101101001010 : data = 16'b1111110000101100;
            15'b000101101001011 : data = 16'b1111110000100111;
            15'b000101101001100 : data = 16'b1111110000100010;
            15'b000101101001101 : data = 16'b1111110000011101;
            15'b000101101001110 : data = 16'b1111110000011000;
            15'b000101101001111 : data = 16'b1111110000010011;
            15'b000101101010000 : data = 16'b1111110000001101;
            15'b000101101010001 : data = 16'b1111110000001000;
            15'b000101101010010 : data = 16'b1111110000000011;
            15'b000101101010011 : data = 16'b1111101111111110;
            15'b000101101010100 : data = 16'b1111101111111001;
            15'b000101101010101 : data = 16'b1111101111110100;
            15'b000101101010110 : data = 16'b1111101111101111;
            15'b000101101010111 : data = 16'b1111101111101010;
            15'b000101101011000 : data = 16'b1111101111100100;
            15'b000101101011001 : data = 16'b1111101111011111;
            15'b000101101011010 : data = 16'b1111101111011010;
            15'b000101101011011 : data = 16'b1111101111010101;
            15'b000101101011100 : data = 16'b1111101111010000;
            15'b000101101011101 : data = 16'b1111101111001010;
            15'b000101101011110 : data = 16'b1111101111000101;
            15'b000101101011111 : data = 16'b1111101111000000;
            15'b000101101100000 : data = 16'b1111101110111011;
            15'b000101101100001 : data = 16'b1111101110110101;
            15'b000101101100010 : data = 16'b1111101110110000;
            15'b000101101100011 : data = 16'b1111101110101011;
            15'b000101101100100 : data = 16'b1111101110100110;
            15'b000101101100101 : data = 16'b1111101110100000;
            15'b000101101100110 : data = 16'b1111101110011011;
            15'b000101101100111 : data = 16'b1111101110010110;
            15'b000101101101000 : data = 16'b1111101110010000;
            15'b000101101101001 : data = 16'b1111101110001011;
            15'b000101101101010 : data = 16'b1111101110000101;
            15'b000101101101011 : data = 16'b1111101110000000;
            15'b000101101101100 : data = 16'b1111101101111011;
            15'b000101101101101 : data = 16'b1111101101110101;
            15'b000101101101110 : data = 16'b1111101101110000;
            15'b000101101101111 : data = 16'b1111101101101010;
            15'b000101101110000 : data = 16'b1111101101100101;
            15'b000101101110001 : data = 16'b1111101101011111;
            15'b000101101110010 : data = 16'b1111101101011010;
            15'b000101101110011 : data = 16'b1111101101010100;
            15'b000101101110100 : data = 16'b1111101101001111;
            15'b000101101110101 : data = 16'b1111101101001001;
            15'b000101101110110 : data = 16'b1111101101000100;
            15'b000101101110111 : data = 16'b1111101100111110;
            15'b000101101111000 : data = 16'b1111101100111001;
            15'b000101101111001 : data = 16'b1111101100110011;
            15'b000101101111010 : data = 16'b1111101100101101;
            15'b000101101111011 : data = 16'b1111101100101000;
            15'b000101101111100 : data = 16'b1111101100100010;
            15'b000101101111101 : data = 16'b1111101100011101;
            15'b000101101111110 : data = 16'b1111101100010111;
            15'b000101101111111 : data = 16'b1111101100010001;
            15'b000101110000000 : data = 16'b1111101100001100;
            15'b000101110000001 : data = 16'b1111101100000110;
            15'b000101110000010 : data = 16'b1111101100000000;
            15'b000101110000011 : data = 16'b1111101011111011;
            15'b000101110000100 : data = 16'b1111101011110101;
            15'b000101110000101 : data = 16'b1111101011101111;
            15'b000101110000110 : data = 16'b1111101011101001;
            15'b000101110000111 : data = 16'b1111101011100100;
            15'b000101110001000 : data = 16'b1111101011011110;
            15'b000101110001001 : data = 16'b1111101011011000;
            15'b000101110001010 : data = 16'b1111101011010010;
            15'b000101110001011 : data = 16'b1111101011001101;
            15'b000101110001100 : data = 16'b1111101011000111;
            15'b000101110001101 : data = 16'b1111101011000001;
            15'b000101110001110 : data = 16'b1111101010111011;
            15'b000101110001111 : data = 16'b1111101010110101;
            15'b000101110010000 : data = 16'b1111101010101111;
            15'b000101110010001 : data = 16'b1111101010101010;
            15'b000101110010010 : data = 16'b1111101010100100;
            15'b000101110010011 : data = 16'b1111101010011110;
            15'b000101110010100 : data = 16'b1111101010011000;
            15'b000101110010101 : data = 16'b1111101010010010;
            15'b000101110010110 : data = 16'b1111101010001100;
            15'b000101110010111 : data = 16'b1111101010000110;
            15'b000101110011000 : data = 16'b1111101010000000;
            15'b000101110011001 : data = 16'b1111101001111010;
            15'b000101110011010 : data = 16'b1111101001110100;
            15'b000101110011011 : data = 16'b1111101001101110;
            15'b000101110011100 : data = 16'b1111101001101000;
            15'b000101110011101 : data = 16'b1111101001100010;
            15'b000101110011110 : data = 16'b1111101001011100;
            15'b000101110011111 : data = 16'b1111101001010110;
            15'b000101110100000 : data = 16'b1111101001010000;
            15'b000101110100001 : data = 16'b1111101001001010;
            15'b000101110100010 : data = 16'b1111101001000100;
            15'b000101110100011 : data = 16'b1111101000111110;
            15'b000101110100100 : data = 16'b1111101000111000;
            15'b000101110100101 : data = 16'b1111101000110001;
            15'b000101110100110 : data = 16'b1111101000101011;
            15'b000101110100111 : data = 16'b1111101000100101;
            15'b000101110101000 : data = 16'b1111101000011111;
            15'b000101110101001 : data = 16'b1111101000011001;
            15'b000101110101010 : data = 16'b1111101000010011;
            15'b000101110101011 : data = 16'b1111101000001100;
            15'b000101110101100 : data = 16'b1111101000000110;
            15'b000101110101101 : data = 16'b1111101000000000;
            15'b000101110101110 : data = 16'b1111100111111010;
            15'b000101110101111 : data = 16'b1111100111110100;
            15'b000101110110000 : data = 16'b1111100111101101;
            15'b000101110110001 : data = 16'b1111100111100111;
            15'b000101110110010 : data = 16'b1111100111100001;
            15'b000101110110011 : data = 16'b1111100111011010;
            15'b000101110110100 : data = 16'b1111100111010100;
            15'b000101110110101 : data = 16'b1111100111001110;
            15'b000101110110110 : data = 16'b1111100111000111;
            15'b000101110110111 : data = 16'b1111100111000001;
            15'b000101110111000 : data = 16'b1111100110111011;
            15'b000101110111001 : data = 16'b1111100110110100;
            15'b000101110111010 : data = 16'b1111100110101110;
            15'b000101110111011 : data = 16'b1111100110101000;
            15'b000101110111100 : data = 16'b1111100110100001;
            15'b000101110111101 : data = 16'b1111100110011011;
            15'b000101110111110 : data = 16'b1111100110010100;
            15'b000101110111111 : data = 16'b1111100110001110;
            15'b000101111000000 : data = 16'b1111100110000111;
            15'b000101111000001 : data = 16'b1111100110000001;
            15'b000101111000010 : data = 16'b1111100101111011;
            15'b000101111000011 : data = 16'b1111100101110100;
            15'b000101111000100 : data = 16'b1111100101101110;
            15'b000101111000101 : data = 16'b1111100101100111;
            15'b000101111000110 : data = 16'b1111100101100000;
            15'b000101111000111 : data = 16'b1111100101011010;
            15'b000101111001000 : data = 16'b1111100101010011;
            15'b000101111001001 : data = 16'b1111100101001101;
            15'b000101111001010 : data = 16'b1111100101000110;
            15'b000101111001011 : data = 16'b1111100101000000;
            15'b000101111001100 : data = 16'b1111100100111001;
            15'b000101111001101 : data = 16'b1111100100110010;
            15'b000101111001110 : data = 16'b1111100100101100;
            15'b000101111001111 : data = 16'b1111100100100101;
            15'b000101111010000 : data = 16'b1111100100011111;
            15'b000101111010001 : data = 16'b1111100100011000;
            15'b000101111010010 : data = 16'b1111100100010001;
            15'b000101111010011 : data = 16'b1111100100001011;
            15'b000101111010100 : data = 16'b1111100100000100;
            15'b000101111010101 : data = 16'b1111100011111101;
            15'b000101111010110 : data = 16'b1111100011110110;
            15'b000101111010111 : data = 16'b1111100011110000;
            15'b000101111011000 : data = 16'b1111100011101001;
            15'b000101111011001 : data = 16'b1111100011100010;
            15'b000101111011010 : data = 16'b1111100011011011;
            15'b000101111011011 : data = 16'b1111100011010101;
            15'b000101111011100 : data = 16'b1111100011001110;
            15'b000101111011101 : data = 16'b1111100011000111;
            15'b000101111011110 : data = 16'b1111100011000000;
            15'b000101111011111 : data = 16'b1111100010111001;
            15'b000101111100000 : data = 16'b1111100010110010;
            15'b000101111100001 : data = 16'b1111100010101100;
            15'b000101111100010 : data = 16'b1111100010100101;
            15'b000101111100011 : data = 16'b1111100010011110;
            15'b000101111100100 : data = 16'b1111100010010111;
            15'b000101111100101 : data = 16'b1111100010010000;
            15'b000101111100110 : data = 16'b1111100010001001;
            15'b000101111100111 : data = 16'b1111100010000010;
            15'b000101111101000 : data = 16'b1111100001111011;
            15'b000101111101001 : data = 16'b1111100001110100;
            15'b000101111101010 : data = 16'b1111100001101101;
            15'b000101111101011 : data = 16'b1111100001100110;
            15'b000101111101100 : data = 16'b1111100001011111;
            15'b000101111101101 : data = 16'b1111100001011000;
            15'b000101111101110 : data = 16'b1111100001010001;
            15'b000101111101111 : data = 16'b1111100001001010;
            15'b000101111110000 : data = 16'b1111100001000011;
            15'b000101111110001 : data = 16'b1111100000111100;
            15'b000101111110010 : data = 16'b1111100000110101;
            15'b000101111110011 : data = 16'b1111100000101110;
            15'b000101111110100 : data = 16'b1111100000100111;
            15'b000101111110101 : data = 16'b1111100000100000;
            15'b000101111110110 : data = 16'b1111100000011001;
            15'b000101111110111 : data = 16'b1111100000010010;
            15'b000101111111000 : data = 16'b1111100000001011;
            15'b000101111111001 : data = 16'b1111100000000011;
            15'b000101111111010 : data = 16'b1111011111111100;
            15'b000101111111011 : data = 16'b1111011111110101;
            15'b000101111111100 : data = 16'b1111011111101110;
            15'b000101111111101 : data = 16'b1111011111100111;
            15'b000101111111110 : data = 16'b1111011111011111;
            15'b000101111111111 : data = 16'b1111011111011000;
            15'b000110000000000 : data = 16'b1111011111010001;
            15'b000110000000001 : data = 16'b1111011111001010;
            15'b000110000000010 : data = 16'b1111011111000010;
            15'b000110000000011 : data = 16'b1111011110111011;
            15'b000110000000100 : data = 16'b1111011110110100;
            15'b000110000000101 : data = 16'b1111011110101101;
            15'b000110000000110 : data = 16'b1111011110100101;
            15'b000110000000111 : data = 16'b1111011110011110;
            15'b000110000001000 : data = 16'b1111011110010111;
            15'b000110000001001 : data = 16'b1111011110001111;
            15'b000110000001010 : data = 16'b1111011110001000;
            15'b000110000001011 : data = 16'b1111011110000001;
            15'b000110000001100 : data = 16'b1111011101111001;
            15'b000110000001101 : data = 16'b1111011101110010;
            15'b000110000001110 : data = 16'b1111011101101010;
            15'b000110000001111 : data = 16'b1111011101100011;
            15'b000110000010000 : data = 16'b1111011101011100;
            15'b000110000010001 : data = 16'b1111011101010100;
            15'b000110000010010 : data = 16'b1111011101001101;
            15'b000110000010011 : data = 16'b1111011101000101;
            15'b000110000010100 : data = 16'b1111011100111110;
            15'b000110000010101 : data = 16'b1111011100110110;
            15'b000110000010110 : data = 16'b1111011100101111;
            15'b000110000010111 : data = 16'b1111011100100111;
            15'b000110000011000 : data = 16'b1111011100100000;
            15'b000110000011001 : data = 16'b1111011100011000;
            15'b000110000011010 : data = 16'b1111011100010001;
            15'b000110000011011 : data = 16'b1111011100001001;
            15'b000110000011100 : data = 16'b1111011100000001;
            15'b000110000011101 : data = 16'b1111011011111010;
            15'b000110000011110 : data = 16'b1111011011110010;
            15'b000110000011111 : data = 16'b1111011011101011;
            15'b000110000100000 : data = 16'b1111011011100011;
            15'b000110000100001 : data = 16'b1111011011011011;
            15'b000110000100010 : data = 16'b1111011011010100;
            15'b000110000100011 : data = 16'b1111011011001100;
            15'b000110000100100 : data = 16'b1111011011000100;
            15'b000110000100101 : data = 16'b1111011010111101;
            15'b000110000100110 : data = 16'b1111011010110101;
            15'b000110000100111 : data = 16'b1111011010101101;
            15'b000110000101000 : data = 16'b1111011010100110;
            15'b000110000101001 : data = 16'b1111011010011110;
            15'b000110000101010 : data = 16'b1111011010010110;
            15'b000110000101011 : data = 16'b1111011010001110;
            15'b000110000101100 : data = 16'b1111011010000111;
            15'b000110000101101 : data = 16'b1111011001111111;
            15'b000110000101110 : data = 16'b1111011001110111;
            15'b000110000101111 : data = 16'b1111011001101111;
            15'b000110000110000 : data = 16'b1111011001101000;
            15'b000110000110001 : data = 16'b1111011001100000;
            15'b000110000110010 : data = 16'b1111011001011000;
            15'b000110000110011 : data = 16'b1111011001010000;
            15'b000110000110100 : data = 16'b1111011001001000;
            15'b000110000110101 : data = 16'b1111011001000000;
            15'b000110000110110 : data = 16'b1111011000111000;
            15'b000110000110111 : data = 16'b1111011000110000;
            15'b000110000111000 : data = 16'b1111011000101001;
            15'b000110000111001 : data = 16'b1111011000100001;
            15'b000110000111010 : data = 16'b1111011000011001;
            15'b000110000111011 : data = 16'b1111011000010001;
            15'b000110000111100 : data = 16'b1111011000001001;
            15'b000110000111101 : data = 16'b1111011000000001;
            15'b000110000111110 : data = 16'b1111010111111001;
            15'b000110000111111 : data = 16'b1111010111110001;
            15'b000110001000000 : data = 16'b1111010111101001;
            15'b000110001000001 : data = 16'b1111010111100001;
            15'b000110001000010 : data = 16'b1111010111011001;
            15'b000110001000011 : data = 16'b1111010111010001;
            15'b000110001000100 : data = 16'b1111010111001001;
            15'b000110001000101 : data = 16'b1111010111000001;
            15'b000110001000110 : data = 16'b1111010110111001;
            15'b000110001000111 : data = 16'b1111010110110001;
            15'b000110001001000 : data = 16'b1111010110101000;
            15'b000110001001001 : data = 16'b1111010110100000;
            15'b000110001001010 : data = 16'b1111010110011000;
            15'b000110001001011 : data = 16'b1111010110010000;
            15'b000110001001100 : data = 16'b1111010110001000;
            15'b000110001001101 : data = 16'b1111010110000000;
            15'b000110001001110 : data = 16'b1111010101111000;
            15'b000110001001111 : data = 16'b1111010101101111;
            15'b000110001010000 : data = 16'b1111010101100111;
            15'b000110001010001 : data = 16'b1111010101011111;
            15'b000110001010010 : data = 16'b1111010101010111;
            15'b000110001010011 : data = 16'b1111010101001111;
            15'b000110001010100 : data = 16'b1111010101000110;
            15'b000110001010101 : data = 16'b1111010100111110;
            15'b000110001010110 : data = 16'b1111010100110110;
            15'b000110001010111 : data = 16'b1111010100101101;
            15'b000110001011000 : data = 16'b1111010100100101;
            15'b000110001011001 : data = 16'b1111010100011101;
            15'b000110001011010 : data = 16'b1111010100010101;
            15'b000110001011011 : data = 16'b1111010100001100;
            15'b000110001011100 : data = 16'b1111010100000100;
            15'b000110001011101 : data = 16'b1111010011111100;
            15'b000110001011110 : data = 16'b1111010011110011;
            15'b000110001011111 : data = 16'b1111010011101011;
            15'b000110001100000 : data = 16'b1111010011100010;
            15'b000110001100001 : data = 16'b1111010011011010;
            15'b000110001100010 : data = 16'b1111010011010010;
            15'b000110001100011 : data = 16'b1111010011001001;
            15'b000110001100100 : data = 16'b1111010011000001;
            15'b000110001100101 : data = 16'b1111010010111000;
            15'b000110001100110 : data = 16'b1111010010110000;
            15'b000110001100111 : data = 16'b1111010010100111;
            15'b000110001101000 : data = 16'b1111010010011111;
            15'b000110001101001 : data = 16'b1111010010010110;
            15'b000110001101010 : data = 16'b1111010010001110;
            15'b000110001101011 : data = 16'b1111010010000101;
            15'b000110001101100 : data = 16'b1111010001111101;
            15'b000110001101101 : data = 16'b1111010001110100;
            15'b000110001101110 : data = 16'b1111010001101100;
            15'b000110001101111 : data = 16'b1111010001100011;
            15'b000110001110000 : data = 16'b1111010001011011;
            15'b000110001110001 : data = 16'b1111010001010010;
            15'b000110001110010 : data = 16'b1111010001001010;
            15'b000110001110011 : data = 16'b1111010001000001;
            15'b000110001110100 : data = 16'b1111010000111000;
            15'b000110001110101 : data = 16'b1111010000110000;
            15'b000110001110110 : data = 16'b1111010000100111;
            15'b000110001110111 : data = 16'b1111010000011110;
            15'b000110001111000 : data = 16'b1111010000010110;
            15'b000110001111001 : data = 16'b1111010000001101;
            15'b000110001111010 : data = 16'b1111010000000100;
            15'b000110001111011 : data = 16'b1111001111111100;
            15'b000110001111100 : data = 16'b1111001111110011;
            15'b000110001111101 : data = 16'b1111001111101010;
            15'b000110001111110 : data = 16'b1111001111100001;
            15'b000110001111111 : data = 16'b1111001111011001;
            15'b000110010000000 : data = 16'b1111001111010000;
            15'b000110010000001 : data = 16'b1111001111000111;
            15'b000110010000010 : data = 16'b1111001110111110;
            15'b000110010000011 : data = 16'b1111001110110110;
            15'b000110010000100 : data = 16'b1111001110101101;
            15'b000110010000101 : data = 16'b1111001110100100;
            15'b000110010000110 : data = 16'b1111001110011011;
            15'b000110010000111 : data = 16'b1111001110010010;
            15'b000110010001000 : data = 16'b1111001110001001;
            15'b000110010001001 : data = 16'b1111001110000001;
            15'b000110010001010 : data = 16'b1111001101111000;
            15'b000110010001011 : data = 16'b1111001101101111;
            15'b000110010001100 : data = 16'b1111001101100110;
            15'b000110010001101 : data = 16'b1111001101011101;
            15'b000110010001110 : data = 16'b1111001101010100;
            15'b000110010001111 : data = 16'b1111001101001011;
            15'b000110010010000 : data = 16'b1111001101000010;
            15'b000110010010001 : data = 16'b1111001100111001;
            15'b000110010010010 : data = 16'b1111001100110000;
            15'b000110010010011 : data = 16'b1111001100100111;
            15'b000110010010100 : data = 16'b1111001100011110;
            15'b000110010010101 : data = 16'b1111001100010101;
            15'b000110010010110 : data = 16'b1111001100001100;
            15'b000110010010111 : data = 16'b1111001100000011;
            15'b000110010011000 : data = 16'b1111001011111010;
            15'b000110010011001 : data = 16'b1111001011110001;
            15'b000110010011010 : data = 16'b1111001011101000;
            15'b000110010011011 : data = 16'b1111001011011111;
            15'b000110010011100 : data = 16'b1111001011010110;
            15'b000110010011101 : data = 16'b1111001011001101;
            15'b000110010011110 : data = 16'b1111001011000100;
            15'b000110010011111 : data = 16'b1111001010111011;
            15'b000110010100000 : data = 16'b1111001010110001;
            15'b000110010100001 : data = 16'b1111001010101000;
            15'b000110010100010 : data = 16'b1111001010011111;
            15'b000110010100011 : data = 16'b1111001010010110;
            15'b000110010100100 : data = 16'b1111001010001101;
            15'b000110010100101 : data = 16'b1111001010000100;
            15'b000110010100110 : data = 16'b1111001001111010;
            15'b000110010100111 : data = 16'b1111001001110001;
            15'b000110010101000 : data = 16'b1111001001101000;
            15'b000110010101001 : data = 16'b1111001001011111;
            15'b000110010101010 : data = 16'b1111001001010110;
            15'b000110010101011 : data = 16'b1111001001001100;
            15'b000110010101100 : data = 16'b1111001001000011;
            15'b000110010101101 : data = 16'b1111001000111010;
            15'b000110010101110 : data = 16'b1111001000110000;
            15'b000110010101111 : data = 16'b1111001000100111;
            15'b000110010110000 : data = 16'b1111001000011110;
            15'b000110010110001 : data = 16'b1111001000010100;
            15'b000110010110010 : data = 16'b1111001000001011;
            15'b000110010110011 : data = 16'b1111001000000010;
            15'b000110010110100 : data = 16'b1111000111111000;
            15'b000110010110101 : data = 16'b1111000111101111;
            15'b000110010110110 : data = 16'b1111000111100110;
            15'b000110010110111 : data = 16'b1111000111011100;
            15'b000110010111000 : data = 16'b1111000111010011;
            15'b000110010111001 : data = 16'b1111000111001001;
            15'b000110010111010 : data = 16'b1111000111000000;
            15'b000110010111011 : data = 16'b1111000110110111;
            15'b000110010111100 : data = 16'b1111000110101101;
            15'b000110010111101 : data = 16'b1111000110100100;
            15'b000110010111110 : data = 16'b1111000110011010;
            15'b000110010111111 : data = 16'b1111000110010001;
            15'b000110011000000 : data = 16'b1111000110000111;
            15'b000110011000001 : data = 16'b1111000101111110;
            15'b000110011000010 : data = 16'b1111000101110100;
            15'b000110011000011 : data = 16'b1111000101101011;
            15'b000110011000100 : data = 16'b1111000101100001;
            15'b000110011000101 : data = 16'b1111000101010111;
            15'b000110011000110 : data = 16'b1111000101001110;
            15'b000110011000111 : data = 16'b1111000101000100;
            15'b000110011001000 : data = 16'b1111000100111011;
            15'b000110011001001 : data = 16'b1111000100110001;
            15'b000110011001010 : data = 16'b1111000100100111;
            15'b000110011001011 : data = 16'b1111000100011110;
            15'b000110011001100 : data = 16'b1111000100010100;
            15'b000110011001101 : data = 16'b1111000100001011;
            15'b000110011001110 : data = 16'b1111000100000001;
            15'b000110011001111 : data = 16'b1111000011110111;
            15'b000110011010000 : data = 16'b1111000011101110;
            15'b000110011010001 : data = 16'b1111000011100100;
            15'b000110011010010 : data = 16'b1111000011011010;
            15'b000110011010011 : data = 16'b1111000011010000;
            15'b000110011010100 : data = 16'b1111000011000111;
            15'b000110011010101 : data = 16'b1111000010111101;
            15'b000110011010110 : data = 16'b1111000010110011;
            15'b000110011010111 : data = 16'b1111000010101001;
            15'b000110011011000 : data = 16'b1111000010100000;
            15'b000110011011001 : data = 16'b1111000010010110;
            15'b000110011011010 : data = 16'b1111000010001100;
            15'b000110011011011 : data = 16'b1111000010000010;
            15'b000110011011100 : data = 16'b1111000001111000;
            15'b000110011011101 : data = 16'b1111000001101111;
            15'b000110011011110 : data = 16'b1111000001100101;
            15'b000110011011111 : data = 16'b1111000001011011;
            15'b000110011100000 : data = 16'b1111000001010001;
            15'b000110011100001 : data = 16'b1111000001000111;
            15'b000110011100010 : data = 16'b1111000000111101;
            15'b000110011100011 : data = 16'b1111000000110011;
            15'b000110011100100 : data = 16'b1111000000101001;
            15'b000110011100101 : data = 16'b1111000000100000;
            15'b000110011100110 : data = 16'b1111000000010110;
            15'b000110011100111 : data = 16'b1111000000001100;
            15'b000110011101000 : data = 16'b1111000000000010;
            15'b000110011101001 : data = 16'b1110111111111000;
            15'b000110011101010 : data = 16'b1110111111101110;
            15'b000110011101011 : data = 16'b1110111111100100;
            15'b000110011101100 : data = 16'b1110111111011010;
            15'b000110011101101 : data = 16'b1110111111010000;
            15'b000110011101110 : data = 16'b1110111111000110;
            15'b000110011101111 : data = 16'b1110111110111100;
            15'b000110011110000 : data = 16'b1110111110110010;
            15'b000110011110001 : data = 16'b1110111110101000;
            15'b000110011110010 : data = 16'b1110111110011101;
            15'b000110011110011 : data = 16'b1110111110010011;
            15'b000110011110100 : data = 16'b1110111110001001;
            15'b000110011110101 : data = 16'b1110111101111111;
            15'b000110011110110 : data = 16'b1110111101110101;
            15'b000110011110111 : data = 16'b1110111101101011;
            15'b000110011111000 : data = 16'b1110111101100001;
            15'b000110011111001 : data = 16'b1110111101010111;
            15'b000110011111010 : data = 16'b1110111101001100;
            15'b000110011111011 : data = 16'b1110111101000010;
            15'b000110011111100 : data = 16'b1110111100111000;
            15'b000110011111101 : data = 16'b1110111100101110;
            15'b000110011111110 : data = 16'b1110111100100100;
            15'b000110011111111 : data = 16'b1110111100011010;
            15'b000110100000000 : data = 16'b1110111100001111;
            15'b000110100000001 : data = 16'b1110111100000101;
            15'b000110100000010 : data = 16'b1110111011111011;
            15'b000110100000011 : data = 16'b1110111011110001;
            15'b000110100000100 : data = 16'b1110111011100110;
            15'b000110100000101 : data = 16'b1110111011011100;
            15'b000110100000110 : data = 16'b1110111011010010;
            15'b000110100000111 : data = 16'b1110111011000111;
            15'b000110100001000 : data = 16'b1110111010111101;
            15'b000110100001001 : data = 16'b1110111010110011;
            15'b000110100001010 : data = 16'b1110111010101000;
            15'b000110100001011 : data = 16'b1110111010011110;
            15'b000110100001100 : data = 16'b1110111010010100;
            15'b000110100001101 : data = 16'b1110111010001001;
            15'b000110100001110 : data = 16'b1110111001111111;
            15'b000110100001111 : data = 16'b1110111001110101;
            15'b000110100010000 : data = 16'b1110111001101010;
            15'b000110100010001 : data = 16'b1110111001100000;
            15'b000110100010010 : data = 16'b1110111001010101;
            15'b000110100010011 : data = 16'b1110111001001011;
            15'b000110100010100 : data = 16'b1110111001000000;
            15'b000110100010101 : data = 16'b1110111000110110;
            15'b000110100010110 : data = 16'b1110111000101011;
            15'b000110100010111 : data = 16'b1110111000100001;
            15'b000110100011000 : data = 16'b1110111000010110;
            15'b000110100011001 : data = 16'b1110111000001100;
            15'b000110100011010 : data = 16'b1110111000000001;
            15'b000110100011011 : data = 16'b1110110111110111;
            15'b000110100011100 : data = 16'b1110110111101100;
            15'b000110100011101 : data = 16'b1110110111100010;
            15'b000110100011110 : data = 16'b1110110111010111;
            15'b000110100011111 : data = 16'b1110110111001101;
            15'b000110100100000 : data = 16'b1110110111000010;
            15'b000110100100001 : data = 16'b1110110110110111;
            15'b000110100100010 : data = 16'b1110110110101101;
            15'b000110100100011 : data = 16'b1110110110100010;
            15'b000110100100100 : data = 16'b1110110110011000;
            15'b000110100100101 : data = 16'b1110110110001101;
            15'b000110100100110 : data = 16'b1110110110000010;
            15'b000110100100111 : data = 16'b1110110101111000;
            15'b000110100101000 : data = 16'b1110110101101101;
            15'b000110100101001 : data = 16'b1110110101100010;
            15'b000110100101010 : data = 16'b1110110101011000;
            15'b000110100101011 : data = 16'b1110110101001101;
            15'b000110100101100 : data = 16'b1110110101000010;
            15'b000110100101101 : data = 16'b1110110100110111;
            15'b000110100101110 : data = 16'b1110110100101101;
            15'b000110100101111 : data = 16'b1110110100100010;
            15'b000110100110000 : data = 16'b1110110100010111;
            15'b000110100110001 : data = 16'b1110110100001100;
            15'b000110100110010 : data = 16'b1110110100000010;
            15'b000110100110011 : data = 16'b1110110011110111;
            15'b000110100110100 : data = 16'b1110110011101100;
            15'b000110100110101 : data = 16'b1110110011100001;
            15'b000110100110110 : data = 16'b1110110011010110;
            15'b000110100110111 : data = 16'b1110110011001100;
            15'b000110100111000 : data = 16'b1110110011000001;
            15'b000110100111001 : data = 16'b1110110010110110;
            15'b000110100111010 : data = 16'b1110110010101011;
            15'b000110100111011 : data = 16'b1110110010100000;
            15'b000110100111100 : data = 16'b1110110010010101;
            15'b000110100111101 : data = 16'b1110110010001010;
            15'b000110100111110 : data = 16'b1110110001111111;
            15'b000110100111111 : data = 16'b1110110001110100;
            15'b000110101000000 : data = 16'b1110110001101001;
            15'b000110101000001 : data = 16'b1110110001011111;
            15'b000110101000010 : data = 16'b1110110001010100;
            15'b000110101000011 : data = 16'b1110110001001001;
            15'b000110101000100 : data = 16'b1110110000111110;
            15'b000110101000101 : data = 16'b1110110000110011;
            15'b000110101000110 : data = 16'b1110110000101000;
            15'b000110101000111 : data = 16'b1110110000011101;
            15'b000110101001000 : data = 16'b1110110000010010;
            15'b000110101001001 : data = 16'b1110110000000111;
            15'b000110101001010 : data = 16'b1110101111111100;
            15'b000110101001011 : data = 16'b1110101111110000;
            15'b000110101001100 : data = 16'b1110101111100101;
            15'b000110101001101 : data = 16'b1110101111011010;
            15'b000110101001110 : data = 16'b1110101111001111;
            15'b000110101001111 : data = 16'b1110101111000100;
            15'b000110101010000 : data = 16'b1110101110111001;
            15'b000110101010001 : data = 16'b1110101110101110;
            15'b000110101010010 : data = 16'b1110101110100011;
            15'b000110101010011 : data = 16'b1110101110011000;
            15'b000110101010100 : data = 16'b1110101110001100;
            15'b000110101010101 : data = 16'b1110101110000001;
            15'b000110101010110 : data = 16'b1110101101110110;
            15'b000110101010111 : data = 16'b1110101101101011;
            15'b000110101011000 : data = 16'b1110101101100000;
            15'b000110101011001 : data = 16'b1110101101010100;
            15'b000110101011010 : data = 16'b1110101101001001;
            15'b000110101011011 : data = 16'b1110101100111110;
            15'b000110101011100 : data = 16'b1110101100110011;
            15'b000110101011101 : data = 16'b1110101100101000;
            15'b000110101011110 : data = 16'b1110101100011100;
            15'b000110101011111 : data = 16'b1110101100010001;
            15'b000110101100000 : data = 16'b1110101100000110;
            15'b000110101100001 : data = 16'b1110101011111010;
            15'b000110101100010 : data = 16'b1110101011101111;
            15'b000110101100011 : data = 16'b1110101011100100;
            15'b000110101100100 : data = 16'b1110101011011000;
            15'b000110101100101 : data = 16'b1110101011001101;
            15'b000110101100110 : data = 16'b1110101011000010;
            15'b000110101100111 : data = 16'b1110101010110110;
            15'b000110101101000 : data = 16'b1110101010101011;
            15'b000110101101001 : data = 16'b1110101010100000;
            15'b000110101101010 : data = 16'b1110101010010100;
            15'b000110101101011 : data = 16'b1110101010001001;
            15'b000110101101100 : data = 16'b1110101001111101;
            15'b000110101101101 : data = 16'b1110101001110010;
            15'b000110101101110 : data = 16'b1110101001100111;
            15'b000110101101111 : data = 16'b1110101001011011;
            15'b000110101110000 : data = 16'b1110101001010000;
            15'b000110101110001 : data = 16'b1110101001000100;
            15'b000110101110010 : data = 16'b1110101000111001;
            15'b000110101110011 : data = 16'b1110101000101101;
            15'b000110101110100 : data = 16'b1110101000100010;
            15'b000110101110101 : data = 16'b1110101000010110;
            15'b000110101110110 : data = 16'b1110101000001011;
            15'b000110101110111 : data = 16'b1110100111111111;
            15'b000110101111000 : data = 16'b1110100111110100;
            15'b000110101111001 : data = 16'b1110100111101000;
            15'b000110101111010 : data = 16'b1110100111011100;
            15'b000110101111011 : data = 16'b1110100111010001;
            15'b000110101111100 : data = 16'b1110100111000101;
            15'b000110101111101 : data = 16'b1110100110111010;
            15'b000110101111110 : data = 16'b1110100110101110;
            15'b000110101111111 : data = 16'b1110100110100010;
            15'b000110110000000 : data = 16'b1110100110010111;
            15'b000110110000001 : data = 16'b1110100110001011;
            15'b000110110000010 : data = 16'b1110100110000000;
            15'b000110110000011 : data = 16'b1110100101110100;
            15'b000110110000100 : data = 16'b1110100101101000;
            15'b000110110000101 : data = 16'b1110100101011101;
            15'b000110110000110 : data = 16'b1110100101010001;
            15'b000110110000111 : data = 16'b1110100101000101;
            15'b000110110001000 : data = 16'b1110100100111001;
            15'b000110110001001 : data = 16'b1110100100101110;
            15'b000110110001010 : data = 16'b1110100100100010;
            15'b000110110001011 : data = 16'b1110100100010110;
            15'b000110110001100 : data = 16'b1110100100001010;
            15'b000110110001101 : data = 16'b1110100011111111;
            15'b000110110001110 : data = 16'b1110100011110011;
            15'b000110110001111 : data = 16'b1110100011100111;
            15'b000110110010000 : data = 16'b1110100011011011;
            15'b000110110010001 : data = 16'b1110100011001111;
            15'b000110110010010 : data = 16'b1110100011000100;
            15'b000110110010011 : data = 16'b1110100010111000;
            15'b000110110010100 : data = 16'b1110100010101100;
            15'b000110110010101 : data = 16'b1110100010100000;
            15'b000110110010110 : data = 16'b1110100010010100;
            15'b000110110010111 : data = 16'b1110100010001000;
            15'b000110110011000 : data = 16'b1110100001111100;
            15'b000110110011001 : data = 16'b1110100001110001;
            15'b000110110011010 : data = 16'b1110100001100101;
            15'b000110110011011 : data = 16'b1110100001011001;
            15'b000110110011100 : data = 16'b1110100001001101;
            15'b000110110011101 : data = 16'b1110100001000001;
            15'b000110110011110 : data = 16'b1110100000110101;
            15'b000110110011111 : data = 16'b1110100000101001;
            15'b000110110100000 : data = 16'b1110100000011101;
            15'b000110110100001 : data = 16'b1110100000010001;
            15'b000110110100010 : data = 16'b1110100000000101;
            15'b000110110100011 : data = 16'b1110011111111001;
            15'b000110110100100 : data = 16'b1110011111101101;
            15'b000110110100101 : data = 16'b1110011111100001;
            15'b000110110100110 : data = 16'b1110011111010101;
            15'b000110110100111 : data = 16'b1110011111001001;
            15'b000110110101000 : data = 16'b1110011110111101;
            15'b000110110101001 : data = 16'b1110011110110001;
            15'b000110110101010 : data = 16'b1110011110100101;
            15'b000110110101011 : data = 16'b1110011110011001;
            15'b000110110101100 : data = 16'b1110011110001101;
            15'b000110110101101 : data = 16'b1110011110000000;
            15'b000110110101110 : data = 16'b1110011101110100;
            15'b000110110101111 : data = 16'b1110011101101000;
            15'b000110110110000 : data = 16'b1110011101011100;
            15'b000110110110001 : data = 16'b1110011101010000;
            15'b000110110110010 : data = 16'b1110011101000100;
            15'b000110110110011 : data = 16'b1110011100111000;
            15'b000110110110100 : data = 16'b1110011100101011;
            15'b000110110110101 : data = 16'b1110011100011111;
            15'b000110110110110 : data = 16'b1110011100010011;
            15'b000110110110111 : data = 16'b1110011100000111;
            15'b000110110111000 : data = 16'b1110011011111011;
            15'b000110110111001 : data = 16'b1110011011101110;
            15'b000110110111010 : data = 16'b1110011011100010;
            15'b000110110111011 : data = 16'b1110011011010110;
            15'b000110110111100 : data = 16'b1110011011001010;
            15'b000110110111101 : data = 16'b1110011010111101;
            15'b000110110111110 : data = 16'b1110011010110001;
            15'b000110110111111 : data = 16'b1110011010100101;
            15'b000110111000000 : data = 16'b1110011010011000;
            15'b000110111000001 : data = 16'b1110011010001100;
            15'b000110111000010 : data = 16'b1110011010000000;
            15'b000110111000011 : data = 16'b1110011001110011;
            15'b000110111000100 : data = 16'b1110011001100111;
            15'b000110111000101 : data = 16'b1110011001011011;
            15'b000110111000110 : data = 16'b1110011001001110;
            15'b000110111000111 : data = 16'b1110011001000010;
            15'b000110111001000 : data = 16'b1110011000110110;
            15'b000110111001001 : data = 16'b1110011000101001;
            15'b000110111001010 : data = 16'b1110011000011101;
            15'b000110111001011 : data = 16'b1110011000010000;
            15'b000110111001100 : data = 16'b1110011000000100;
            15'b000110111001101 : data = 16'b1110010111111000;
            15'b000110111001110 : data = 16'b1110010111101011;
            15'b000110111001111 : data = 16'b1110010111011111;
            15'b000110111010000 : data = 16'b1110010111010010;
            15'b000110111010001 : data = 16'b1110010111000110;
            15'b000110111010010 : data = 16'b1110010110111001;
            15'b000110111010011 : data = 16'b1110010110101101;
            15'b000110111010100 : data = 16'b1110010110100000;
            15'b000110111010101 : data = 16'b1110010110010100;
            15'b000110111010110 : data = 16'b1110010110000111;
            15'b000110111010111 : data = 16'b1110010101111011;
            15'b000110111011000 : data = 16'b1110010101101110;
            15'b000110111011001 : data = 16'b1110010101100001;
            15'b000110111011010 : data = 16'b1110010101010101;
            15'b000110111011011 : data = 16'b1110010101001000;
            15'b000110111011100 : data = 16'b1110010100111100;
            15'b000110111011101 : data = 16'b1110010100101111;
            15'b000110111011110 : data = 16'b1110010100100011;
            15'b000110111011111 : data = 16'b1110010100010110;
            15'b000110111100000 : data = 16'b1110010100001001;
            15'b000110111100001 : data = 16'b1110010011111101;
            15'b000110111100010 : data = 16'b1110010011110000;
            15'b000110111100011 : data = 16'b1110010011100011;
            15'b000110111100100 : data = 16'b1110010011010111;
            15'b000110111100101 : data = 16'b1110010011001010;
            15'b000110111100110 : data = 16'b1110010010111101;
            15'b000110111100111 : data = 16'b1110010010110001;
            15'b000110111101000 : data = 16'b1110010010100100;
            15'b000110111101001 : data = 16'b1110010010010111;
            15'b000110111101010 : data = 16'b1110010010001010;
            15'b000110111101011 : data = 16'b1110010001111110;
            15'b000110111101100 : data = 16'b1110010001110001;
            15'b000110111101101 : data = 16'b1110010001100100;
            15'b000110111101110 : data = 16'b1110010001010111;
            15'b000110111101111 : data = 16'b1110010001001011;
            15'b000110111110000 : data = 16'b1110010000111110;
            15'b000110111110001 : data = 16'b1110010000110001;
            15'b000110111110010 : data = 16'b1110010000100100;
            15'b000110111110011 : data = 16'b1110010000010111;
            15'b000110111110100 : data = 16'b1110010000001010;
            15'b000110111110101 : data = 16'b1110001111111110;
            15'b000110111110110 : data = 16'b1110001111110001;
            15'b000110111110111 : data = 16'b1110001111100100;
            15'b000110111111000 : data = 16'b1110001111010111;
            15'b000110111111001 : data = 16'b1110001111001010;
            15'b000110111111010 : data = 16'b1110001110111101;
            15'b000110111111011 : data = 16'b1110001110110000;
            15'b000110111111100 : data = 16'b1110001110100011;
            15'b000110111111101 : data = 16'b1110001110010110;
            15'b000110111111110 : data = 16'b1110001110001010;
            15'b000110111111111 : data = 16'b1110001101111101;
            15'b000111000000000 : data = 16'b1110001101110000;
            15'b000111000000001 : data = 16'b1110001101100011;
            15'b000111000000010 : data = 16'b1110001101010110;
            15'b000111000000011 : data = 16'b1110001101001001;
            15'b000111000000100 : data = 16'b1110001100111100;
            15'b000111000000101 : data = 16'b1110001100101111;
            15'b000111000000110 : data = 16'b1110001100100010;
            15'b000111000000111 : data = 16'b1110001100010101;
            15'b000111000001000 : data = 16'b1110001100001000;
            15'b000111000001001 : data = 16'b1110001011111011;
            15'b000111000001010 : data = 16'b1110001011101101;
            15'b000111000001011 : data = 16'b1110001011100000;
            15'b000111000001100 : data = 16'b1110001011010011;
            15'b000111000001101 : data = 16'b1110001011000110;
            15'b000111000001110 : data = 16'b1110001010111001;
            15'b000111000001111 : data = 16'b1110001010101100;
            15'b000111000010000 : data = 16'b1110001010011111;
            15'b000111000010001 : data = 16'b1110001010010010;
            15'b000111000010010 : data = 16'b1110001010000101;
            15'b000111000010011 : data = 16'b1110001001110111;
            15'b000111000010100 : data = 16'b1110001001101010;
            15'b000111000010101 : data = 16'b1110001001011101;
            15'b000111000010110 : data = 16'b1110001001010000;
            15'b000111000010111 : data = 16'b1110001001000011;
            15'b000111000011000 : data = 16'b1110001000110110;
            15'b000111000011001 : data = 16'b1110001000101000;
            15'b000111000011010 : data = 16'b1110001000011011;
            15'b000111000011011 : data = 16'b1110001000001110;
            15'b000111000011100 : data = 16'b1110001000000001;
            15'b000111000011101 : data = 16'b1110000111110011;
            15'b000111000011110 : data = 16'b1110000111100110;
            15'b000111000011111 : data = 16'b1110000111011001;
            15'b000111000100000 : data = 16'b1110000111001100;
            15'b000111000100001 : data = 16'b1110000110111110;
            15'b000111000100010 : data = 16'b1110000110110001;
            15'b000111000100011 : data = 16'b1110000110100100;
            15'b000111000100100 : data = 16'b1110000110010110;
            15'b000111000100101 : data = 16'b1110000110001001;
            15'b000111000100110 : data = 16'b1110000101111100;
            15'b000111000100111 : data = 16'b1110000101101110;
            15'b000111000101000 : data = 16'b1110000101100001;
            15'b000111000101001 : data = 16'b1110000101010100;
            15'b000111000101010 : data = 16'b1110000101000110;
            15'b000111000101011 : data = 16'b1110000100111001;
            15'b000111000101100 : data = 16'b1110000100101100;
            15'b000111000101101 : data = 16'b1110000100011110;
            15'b000111000101110 : data = 16'b1110000100010001;
            15'b000111000101111 : data = 16'b1110000100000011;
            15'b000111000110000 : data = 16'b1110000011110110;
            15'b000111000110001 : data = 16'b1110000011101000;
            15'b000111000110010 : data = 16'b1110000011011011;
            15'b000111000110011 : data = 16'b1110000011001110;
            15'b000111000110100 : data = 16'b1110000011000000;
            15'b000111000110101 : data = 16'b1110000010110011;
            15'b000111000110110 : data = 16'b1110000010100101;
            15'b000111000110111 : data = 16'b1110000010011000;
            15'b000111000111000 : data = 16'b1110000010001010;
            15'b000111000111001 : data = 16'b1110000001111101;
            15'b000111000111010 : data = 16'b1110000001101111;
            15'b000111000111011 : data = 16'b1110000001100001;
            15'b000111000111100 : data = 16'b1110000001010100;
            15'b000111000111101 : data = 16'b1110000001000110;
            15'b000111000111110 : data = 16'b1110000000111001;
            15'b000111000111111 : data = 16'b1110000000101011;
            15'b000111001000000 : data = 16'b1110000000011110;
            15'b000111001000001 : data = 16'b1110000000010000;
            15'b000111001000010 : data = 16'b1110000000000010;
            15'b000111001000011 : data = 16'b1101111111110101;
            15'b000111001000100 : data = 16'b1101111111100111;
            15'b000111001000101 : data = 16'b1101111111011010;
            15'b000111001000110 : data = 16'b1101111111001100;
            15'b000111001000111 : data = 16'b1101111110111110;
            15'b000111001001000 : data = 16'b1101111110110001;
            15'b000111001001001 : data = 16'b1101111110100011;
            15'b000111001001010 : data = 16'b1101111110010101;
            15'b000111001001011 : data = 16'b1101111110000111;
            15'b000111001001100 : data = 16'b1101111101111010;
            15'b000111001001101 : data = 16'b1101111101101100;
            15'b000111001001110 : data = 16'b1101111101011110;
            15'b000111001001111 : data = 16'b1101111101010001;
            15'b000111001010000 : data = 16'b1101111101000011;
            15'b000111001010001 : data = 16'b1101111100110101;
            15'b000111001010010 : data = 16'b1101111100100111;
            15'b000111001010011 : data = 16'b1101111100011010;
            15'b000111001010100 : data = 16'b1101111100001100;
            15'b000111001010101 : data = 16'b1101111011111110;
            15'b000111001010110 : data = 16'b1101111011110000;
            15'b000111001010111 : data = 16'b1101111011100010;
            15'b000111001011000 : data = 16'b1101111011010101;
            15'b000111001011001 : data = 16'b1101111011000111;
            15'b000111001011010 : data = 16'b1101111010111001;
            15'b000111001011011 : data = 16'b1101111010101011;
            15'b000111001011100 : data = 16'b1101111010011101;
            15'b000111001011101 : data = 16'b1101111010001111;
            15'b000111001011110 : data = 16'b1101111010000001;
            15'b000111001011111 : data = 16'b1101111001110011;
            15'b000111001100000 : data = 16'b1101111001100110;
            15'b000111001100001 : data = 16'b1101111001011000;
            15'b000111001100010 : data = 16'b1101111001001010;
            15'b000111001100011 : data = 16'b1101111000111100;
            15'b000111001100100 : data = 16'b1101111000101110;
            15'b000111001100101 : data = 16'b1101111000100000;
            15'b000111001100110 : data = 16'b1101111000010010;
            15'b000111001100111 : data = 16'b1101111000000100;
            15'b000111001101000 : data = 16'b1101110111110110;
            15'b000111001101001 : data = 16'b1101110111101000;
            15'b000111001101010 : data = 16'b1101110111011010;
            15'b000111001101011 : data = 16'b1101110111001100;
            15'b000111001101100 : data = 16'b1101110110111110;
            15'b000111001101101 : data = 16'b1101110110110000;
            15'b000111001101110 : data = 16'b1101110110100010;
            15'b000111001101111 : data = 16'b1101110110010100;
            15'b000111001110000 : data = 16'b1101110110000110;
            15'b000111001110001 : data = 16'b1101110101111000;
            15'b000111001110010 : data = 16'b1101110101101010;
            15'b000111001110011 : data = 16'b1101110101011100;
            15'b000111001110100 : data = 16'b1101110101001110;
            15'b000111001110101 : data = 16'b1101110101000000;
            15'b000111001110110 : data = 16'b1101110100110001;
            15'b000111001110111 : data = 16'b1101110100100011;
            15'b000111001111000 : data = 16'b1101110100010101;
            15'b000111001111001 : data = 16'b1101110100000111;
            15'b000111001111010 : data = 16'b1101110011111001;
            15'b000111001111011 : data = 16'b1101110011101011;
            15'b000111001111100 : data = 16'b1101110011011101;
            15'b000111001111101 : data = 16'b1101110011001110;
            15'b000111001111110 : data = 16'b1101110011000000;
            15'b000111001111111 : data = 16'b1101110010110010;
            15'b000111010000000 : data = 16'b1101110010100100;
            15'b000111010000001 : data = 16'b1101110010010110;
            15'b000111010000010 : data = 16'b1101110010000111;
            15'b000111010000011 : data = 16'b1101110001111001;
            15'b000111010000100 : data = 16'b1101110001101011;
            15'b000111010000101 : data = 16'b1101110001011101;
            15'b000111010000110 : data = 16'b1101110001001110;
            15'b000111010000111 : data = 16'b1101110001000000;
            15'b000111010001000 : data = 16'b1101110000110010;
            15'b000111010001001 : data = 16'b1101110000100100;
            15'b000111010001010 : data = 16'b1101110000010101;
            15'b000111010001011 : data = 16'b1101110000000111;
            15'b000111010001100 : data = 16'b1101101111111001;
            15'b000111010001101 : data = 16'b1101101111101010;
            15'b000111010001110 : data = 16'b1101101111011100;
            15'b000111010001111 : data = 16'b1101101111001110;
            15'b000111010010000 : data = 16'b1101101110111111;
            15'b000111010010001 : data = 16'b1101101110110001;
            15'b000111010010010 : data = 16'b1101101110100011;
            15'b000111010010011 : data = 16'b1101101110010100;
            15'b000111010010100 : data = 16'b1101101110000110;
            15'b000111010010101 : data = 16'b1101101101110111;
            15'b000111010010110 : data = 16'b1101101101101001;
            15'b000111010010111 : data = 16'b1101101101011011;
            15'b000111010011000 : data = 16'b1101101101001100;
            15'b000111010011001 : data = 16'b1101101100111110;
            15'b000111010011010 : data = 16'b1101101100101111;
            15'b000111010011011 : data = 16'b1101101100100001;
            15'b000111010011100 : data = 16'b1101101100010010;
            15'b000111010011101 : data = 16'b1101101100000100;
            15'b000111010011110 : data = 16'b1101101011110101;
            15'b000111010011111 : data = 16'b1101101011100111;
            15'b000111010100000 : data = 16'b1101101011011000;
            15'b000111010100001 : data = 16'b1101101011001010;
            15'b000111010100010 : data = 16'b1101101010111011;
            15'b000111010100011 : data = 16'b1101101010101101;
            15'b000111010100100 : data = 16'b1101101010011110;
            15'b000111010100101 : data = 16'b1101101010010000;
            15'b000111010100110 : data = 16'b1101101010000001;
            15'b000111010100111 : data = 16'b1101101001110011;
            15'b000111010101000 : data = 16'b1101101001100100;
            15'b000111010101001 : data = 16'b1101101001010110;
            15'b000111010101010 : data = 16'b1101101001000111;
            15'b000111010101011 : data = 16'b1101101000111000;
            15'b000111010101100 : data = 16'b1101101000101010;
            15'b000111010101101 : data = 16'b1101101000011011;
            15'b000111010101110 : data = 16'b1101101000001101;
            15'b000111010101111 : data = 16'b1101100111111110;
            15'b000111010110000 : data = 16'b1101100111101111;
            15'b000111010110001 : data = 16'b1101100111100001;
            15'b000111010110010 : data = 16'b1101100111010010;
            15'b000111010110011 : data = 16'b1101100111000011;
            15'b000111010110100 : data = 16'b1101100110110101;
            15'b000111010110101 : data = 16'b1101100110100110;
            15'b000111010110110 : data = 16'b1101100110010111;
            15'b000111010110111 : data = 16'b1101100110001000;
            15'b000111010111000 : data = 16'b1101100101111010;
            15'b000111010111001 : data = 16'b1101100101101011;
            15'b000111010111010 : data = 16'b1101100101011100;
            15'b000111010111011 : data = 16'b1101100101001110;
            15'b000111010111100 : data = 16'b1101100100111111;
            15'b000111010111101 : data = 16'b1101100100110000;
            15'b000111010111110 : data = 16'b1101100100100001;
            15'b000111010111111 : data = 16'b1101100100010010;
            15'b000111011000000 : data = 16'b1101100100000100;
            15'b000111011000001 : data = 16'b1101100011110101;
            15'b000111011000010 : data = 16'b1101100011100110;
            15'b000111011000011 : data = 16'b1101100011010111;
            15'b000111011000100 : data = 16'b1101100011001000;
            15'b000111011000101 : data = 16'b1101100010111010;
            15'b000111011000110 : data = 16'b1101100010101011;
            15'b000111011000111 : data = 16'b1101100010011100;
            15'b000111011001000 : data = 16'b1101100010001101;
            15'b000111011001001 : data = 16'b1101100001111110;
            15'b000111011001010 : data = 16'b1101100001101111;
            15'b000111011001011 : data = 16'b1101100001100000;
            15'b000111011001100 : data = 16'b1101100001010010;
            15'b000111011001101 : data = 16'b1101100001000011;
            15'b000111011001110 : data = 16'b1101100000110100;
            15'b000111011001111 : data = 16'b1101100000100101;
            15'b000111011010000 : data = 16'b1101100000010110;
            15'b000111011010001 : data = 16'b1101100000000111;
            15'b000111011010010 : data = 16'b1101011111111000;
            15'b000111011010011 : data = 16'b1101011111101001;
            15'b000111011010100 : data = 16'b1101011111011010;
            15'b000111011010101 : data = 16'b1101011111001011;
            15'b000111011010110 : data = 16'b1101011110111100;
            15'b000111011010111 : data = 16'b1101011110101101;
            15'b000111011011000 : data = 16'b1101011110011110;
            15'b000111011011001 : data = 16'b1101011110001111;
            15'b000111011011010 : data = 16'b1101011110000000;
            15'b000111011011011 : data = 16'b1101011101110001;
            15'b000111011011100 : data = 16'b1101011101100010;
            15'b000111011011101 : data = 16'b1101011101010011;
            15'b000111011011110 : data = 16'b1101011101000100;
            15'b000111011011111 : data = 16'b1101011100110101;
            15'b000111011100000 : data = 16'b1101011100100110;
            15'b000111011100001 : data = 16'b1101011100010111;
            15'b000111011100010 : data = 16'b1101011100001000;
            15'b000111011100011 : data = 16'b1101011011111000;
            15'b000111011100100 : data = 16'b1101011011101001;
            15'b000111011100101 : data = 16'b1101011011011010;
            15'b000111011100110 : data = 16'b1101011011001011;
            15'b000111011100111 : data = 16'b1101011010111100;
            15'b000111011101000 : data = 16'b1101011010101101;
            15'b000111011101001 : data = 16'b1101011010011110;
            15'b000111011101010 : data = 16'b1101011010001110;
            15'b000111011101011 : data = 16'b1101011001111111;
            15'b000111011101100 : data = 16'b1101011001110000;
            15'b000111011101101 : data = 16'b1101011001100001;
            15'b000111011101110 : data = 16'b1101011001010010;
            15'b000111011101111 : data = 16'b1101011001000011;
            15'b000111011110000 : data = 16'b1101011000110011;
            15'b000111011110001 : data = 16'b1101011000100100;
            15'b000111011110010 : data = 16'b1101011000010101;
            15'b000111011110011 : data = 16'b1101011000000110;
            15'b000111011110100 : data = 16'b1101010111110110;
            15'b000111011110101 : data = 16'b1101010111100111;
            15'b000111011110110 : data = 16'b1101010111011000;
            15'b000111011110111 : data = 16'b1101010111001001;
            15'b000111011111000 : data = 16'b1101010110111001;
            15'b000111011111001 : data = 16'b1101010110101010;
            15'b000111011111010 : data = 16'b1101010110011011;
            15'b000111011111011 : data = 16'b1101010110001011;
            15'b000111011111100 : data = 16'b1101010101111100;
            15'b000111011111101 : data = 16'b1101010101101101;
            15'b000111011111110 : data = 16'b1101010101011101;
            15'b000111011111111 : data = 16'b1101010101001110;
            15'b000111100000000 : data = 16'b1101010100111111;
            15'b000111100000001 : data = 16'b1101010100101111;
            15'b000111100000010 : data = 16'b1101010100100000;
            15'b000111100000011 : data = 16'b1101010100010001;
            15'b000111100000100 : data = 16'b1101010100000001;
            15'b000111100000101 : data = 16'b1101010011110010;
            15'b000111100000110 : data = 16'b1101010011100010;
            15'b000111100000111 : data = 16'b1101010011010011;
            15'b000111100001000 : data = 16'b1101010011000100;
            15'b000111100001001 : data = 16'b1101010010110100;
            15'b000111100001010 : data = 16'b1101010010100101;
            15'b000111100001011 : data = 16'b1101010010010101;
            15'b000111100001100 : data = 16'b1101010010000110;
            15'b000111100001101 : data = 16'b1101010001110110;
            15'b000111100001110 : data = 16'b1101010001100111;
            15'b000111100001111 : data = 16'b1101010001010111;
            15'b000111100010000 : data = 16'b1101010001001000;
            15'b000111100010001 : data = 16'b1101010000111000;
            15'b000111100010010 : data = 16'b1101010000101001;
            15'b000111100010011 : data = 16'b1101010000011001;
            15'b000111100010100 : data = 16'b1101010000001010;
            15'b000111100010101 : data = 16'b1101001111111010;
            15'b000111100010110 : data = 16'b1101001111101011;
            15'b000111100010111 : data = 16'b1101001111011011;
            15'b000111100011000 : data = 16'b1101001111001100;
            15'b000111100011001 : data = 16'b1101001110111100;
            15'b000111100011010 : data = 16'b1101001110101101;
            15'b000111100011011 : data = 16'b1101001110011101;
            15'b000111100011100 : data = 16'b1101001110001101;
            15'b000111100011101 : data = 16'b1101001101111110;
            15'b000111100011110 : data = 16'b1101001101101110;
            15'b000111100011111 : data = 16'b1101001101011111;
            15'b000111100100000 : data = 16'b1101001101001111;
            15'b000111100100001 : data = 16'b1101001100111111;
            15'b000111100100010 : data = 16'b1101001100110000;
            15'b000111100100011 : data = 16'b1101001100100000;
            15'b000111100100100 : data = 16'b1101001100010000;
            15'b000111100100101 : data = 16'b1101001100000001;
            15'b000111100100110 : data = 16'b1101001011110001;
            15'b000111100100111 : data = 16'b1101001011100001;
            15'b000111100101000 : data = 16'b1101001011010010;
            15'b000111100101001 : data = 16'b1101001011000010;
            15'b000111100101010 : data = 16'b1101001010110010;
            15'b000111100101011 : data = 16'b1101001010100010;
            15'b000111100101100 : data = 16'b1101001010010011;
            15'b000111100101101 : data = 16'b1101001010000011;
            15'b000111100101110 : data = 16'b1101001001110011;
            15'b000111100101111 : data = 16'b1101001001100011;
            15'b000111100110000 : data = 16'b1101001001010100;
            15'b000111100110001 : data = 16'b1101001001000100;
            15'b000111100110010 : data = 16'b1101001000110100;
            15'b000111100110011 : data = 16'b1101001000100100;
            15'b000111100110100 : data = 16'b1101001000010101;
            15'b000111100110101 : data = 16'b1101001000000101;
            15'b000111100110110 : data = 16'b1101000111110101;
            15'b000111100110111 : data = 16'b1101000111100101;
            15'b000111100111000 : data = 16'b1101000111010101;
            15'b000111100111001 : data = 16'b1101000111000110;
            15'b000111100111010 : data = 16'b1101000110110110;
            15'b000111100111011 : data = 16'b1101000110100110;
            15'b000111100111100 : data = 16'b1101000110010110;
            15'b000111100111101 : data = 16'b1101000110000110;
            15'b000111100111110 : data = 16'b1101000101110110;
            15'b000111100111111 : data = 16'b1101000101100110;
            15'b000111101000000 : data = 16'b1101000101010110;
            15'b000111101000001 : data = 16'b1101000101000111;
            15'b000111101000010 : data = 16'b1101000100110111;
            15'b000111101000011 : data = 16'b1101000100100111;
            15'b000111101000100 : data = 16'b1101000100010111;
            15'b000111101000101 : data = 16'b1101000100000111;
            15'b000111101000110 : data = 16'b1101000011110111;
            15'b000111101000111 : data = 16'b1101000011100111;
            15'b000111101001000 : data = 16'b1101000011010111;
            15'b000111101001001 : data = 16'b1101000011000111;
            15'b000111101001010 : data = 16'b1101000010110111;
            15'b000111101001011 : data = 16'b1101000010100111;
            15'b000111101001100 : data = 16'b1101000010010111;
            15'b000111101001101 : data = 16'b1101000010000111;
            15'b000111101001110 : data = 16'b1101000001110111;
            15'b000111101001111 : data = 16'b1101000001100111;
            15'b000111101010000 : data = 16'b1101000001010111;
            15'b000111101010001 : data = 16'b1101000001000111;
            15'b000111101010010 : data = 16'b1101000000110111;
            15'b000111101010011 : data = 16'b1101000000100111;
            15'b000111101010100 : data = 16'b1101000000010111;
            15'b000111101010101 : data = 16'b1101000000000111;
            15'b000111101010110 : data = 16'b1100111111110111;
            15'b000111101010111 : data = 16'b1100111111100111;
            15'b000111101011000 : data = 16'b1100111111010111;
            15'b000111101011001 : data = 16'b1100111111000110;
            15'b000111101011010 : data = 16'b1100111110110110;
            15'b000111101011011 : data = 16'b1100111110100110;
            15'b000111101011100 : data = 16'b1100111110010110;
            15'b000111101011101 : data = 16'b1100111110000110;
            15'b000111101011110 : data = 16'b1100111101110110;
            15'b000111101011111 : data = 16'b1100111101100110;
            15'b000111101100000 : data = 16'b1100111101010110;
            15'b000111101100001 : data = 16'b1100111101000101;
            15'b000111101100010 : data = 16'b1100111100110101;
            15'b000111101100011 : data = 16'b1100111100100101;
            15'b000111101100100 : data = 16'b1100111100010101;
            15'b000111101100101 : data = 16'b1100111100000101;
            15'b000111101100110 : data = 16'b1100111011110101;
            15'b000111101100111 : data = 16'b1100111011100100;
            15'b000111101101000 : data = 16'b1100111011010100;
            15'b000111101101001 : data = 16'b1100111011000100;
            15'b000111101101010 : data = 16'b1100111010110100;
            15'b000111101101011 : data = 16'b1100111010100011;
            15'b000111101101100 : data = 16'b1100111010010011;
            15'b000111101101101 : data = 16'b1100111010000011;
            15'b000111101101110 : data = 16'b1100111001110011;
            15'b000111101101111 : data = 16'b1100111001100010;
            15'b000111101110000 : data = 16'b1100111001010010;
            15'b000111101110001 : data = 16'b1100111001000010;
            15'b000111101110010 : data = 16'b1100111000110001;
            15'b000111101110011 : data = 16'b1100111000100001;
            15'b000111101110100 : data = 16'b1100111000010001;
            15'b000111101110101 : data = 16'b1100111000000001;
            15'b000111101110110 : data = 16'b1100110111110000;
            15'b000111101110111 : data = 16'b1100110111100000;
            15'b000111101111000 : data = 16'b1100110111010000;
            15'b000111101111001 : data = 16'b1100110110111111;
            15'b000111101111010 : data = 16'b1100110110101111;
            15'b000111101111011 : data = 16'b1100110110011110;
            15'b000111101111100 : data = 16'b1100110110001110;
            15'b000111101111101 : data = 16'b1100110101111110;
            15'b000111101111110 : data = 16'b1100110101101101;
            15'b000111101111111 : data = 16'b1100110101011101;
            15'b000111110000000 : data = 16'b1100110101001101;
            15'b000111110000001 : data = 16'b1100110100111100;
            15'b000111110000010 : data = 16'b1100110100101100;
            15'b000111110000011 : data = 16'b1100110100011011;
            15'b000111110000100 : data = 16'b1100110100001011;
            15'b000111110000101 : data = 16'b1100110011111010;
            15'b000111110000110 : data = 16'b1100110011101010;
            15'b000111110000111 : data = 16'b1100110011011001;
            15'b000111110001000 : data = 16'b1100110011001001;
            15'b000111110001001 : data = 16'b1100110010111001;
            15'b000111110001010 : data = 16'b1100110010101000;
            15'b000111110001011 : data = 16'b1100110010011000;
            15'b000111110001100 : data = 16'b1100110010000111;
            15'b000111110001101 : data = 16'b1100110001110111;
            15'b000111110001110 : data = 16'b1100110001100110;
            15'b000111110001111 : data = 16'b1100110001010110;
            15'b000111110010000 : data = 16'b1100110001000101;
            15'b000111110010001 : data = 16'b1100110000110100;
            15'b000111110010010 : data = 16'b1100110000100100;
            15'b000111110010011 : data = 16'b1100110000010011;
            15'b000111110010100 : data = 16'b1100110000000011;
            15'b000111110010101 : data = 16'b1100101111110010;
            15'b000111110010110 : data = 16'b1100101111100010;
            15'b000111110010111 : data = 16'b1100101111010001;
            15'b000111110011000 : data = 16'b1100101111000000;
            15'b000111110011001 : data = 16'b1100101110110000;
            15'b000111110011010 : data = 16'b1100101110011111;
            15'b000111110011011 : data = 16'b1100101110001111;
            15'b000111110011100 : data = 16'b1100101101111110;
            15'b000111110011101 : data = 16'b1100101101101101;
            15'b000111110011110 : data = 16'b1100101101011101;
            15'b000111110011111 : data = 16'b1100101101001100;
            15'b000111110100000 : data = 16'b1100101100111011;
            15'b000111110100001 : data = 16'b1100101100101011;
            15'b000111110100010 : data = 16'b1100101100011010;
            15'b000111110100011 : data = 16'b1100101100001001;
            15'b000111110100100 : data = 16'b1100101011111001;
            15'b000111110100101 : data = 16'b1100101011101000;
            15'b000111110100110 : data = 16'b1100101011010111;
            15'b000111110100111 : data = 16'b1100101011000111;
            15'b000111110101000 : data = 16'b1100101010110110;
            15'b000111110101001 : data = 16'b1100101010100101;
            15'b000111110101010 : data = 16'b1100101010010101;
            15'b000111110101011 : data = 16'b1100101010000100;
            15'b000111110101100 : data = 16'b1100101001110011;
            15'b000111110101101 : data = 16'b1100101001100010;
            15'b000111110101110 : data = 16'b1100101001010010;
            15'b000111110101111 : data = 16'b1100101001000001;
            15'b000111110110000 : data = 16'b1100101000110000;
            15'b000111110110001 : data = 16'b1100101000011111;
            15'b000111110110010 : data = 16'b1100101000001110;
            15'b000111110110011 : data = 16'b1100100111111110;
            15'b000111110110100 : data = 16'b1100100111101101;
            15'b000111110110101 : data = 16'b1100100111011100;
            15'b000111110110110 : data = 16'b1100100111001011;
            15'b000111110110111 : data = 16'b1100100110111010;
            15'b000111110111000 : data = 16'b1100100110101010;
            15'b000111110111001 : data = 16'b1100100110011001;
            15'b000111110111010 : data = 16'b1100100110001000;
            15'b000111110111011 : data = 16'b1100100101110111;
            15'b000111110111100 : data = 16'b1100100101100110;
            15'b000111110111101 : data = 16'b1100100101010101;
            15'b000111110111110 : data = 16'b1100100101000100;
            15'b000111110111111 : data = 16'b1100100100110011;
            15'b000111111000000 : data = 16'b1100100100100011;
            15'b000111111000001 : data = 16'b1100100100010010;
            15'b000111111000010 : data = 16'b1100100100000001;
            15'b000111111000011 : data = 16'b1100100011110000;
            15'b000111111000100 : data = 16'b1100100011011111;
            15'b000111111000101 : data = 16'b1100100011001110;
            15'b000111111000110 : data = 16'b1100100010111101;
            15'b000111111000111 : data = 16'b1100100010101100;
            15'b000111111001000 : data = 16'b1100100010011011;
            15'b000111111001001 : data = 16'b1100100010001010;
            15'b000111111001010 : data = 16'b1100100001111001;
            15'b000111111001011 : data = 16'b1100100001101000;
            15'b000111111001100 : data = 16'b1100100001010111;
            15'b000111111001101 : data = 16'b1100100001000110;
            15'b000111111001110 : data = 16'b1100100000110101;
            15'b000111111001111 : data = 16'b1100100000100100;
            15'b000111111010000 : data = 16'b1100100000010011;
            15'b000111111010001 : data = 16'b1100100000000010;
            15'b000111111010010 : data = 16'b1100011111110001;
            15'b000111111010011 : data = 16'b1100011111100000;
            15'b000111111010100 : data = 16'b1100011111001111;
            15'b000111111010101 : data = 16'b1100011110111110;
            15'b000111111010110 : data = 16'b1100011110101101;
            15'b000111111010111 : data = 16'b1100011110011100;
            15'b000111111011000 : data = 16'b1100011110001011;
            15'b000111111011001 : data = 16'b1100011101111010;
            15'b000111111011010 : data = 16'b1100011101101001;
            15'b000111111011011 : data = 16'b1100011101011000;
            15'b000111111011100 : data = 16'b1100011101000111;
            15'b000111111011101 : data = 16'b1100011100110110;
            15'b000111111011110 : data = 16'b1100011100100100;
            15'b000111111011111 : data = 16'b1100011100010011;
            15'b000111111100000 : data = 16'b1100011100000010;
            15'b000111111100001 : data = 16'b1100011011110001;
            15'b000111111100010 : data = 16'b1100011011100000;
            15'b000111111100011 : data = 16'b1100011011001111;
            15'b000111111100100 : data = 16'b1100011010111110;
            15'b000111111100101 : data = 16'b1100011010101100;
            15'b000111111100110 : data = 16'b1100011010011011;
            15'b000111111100111 : data = 16'b1100011010001010;
            15'b000111111101000 : data = 16'b1100011001111001;
            15'b000111111101001 : data = 16'b1100011001101000;
            15'b000111111101010 : data = 16'b1100011001010111;
            15'b000111111101011 : data = 16'b1100011001000101;
            15'b000111111101100 : data = 16'b1100011000110100;
            15'b000111111101101 : data = 16'b1100011000100011;
            15'b000111111101110 : data = 16'b1100011000010010;
            15'b000111111101111 : data = 16'b1100011000000000;
            15'b000111111110000 : data = 16'b1100010111101111;
            15'b000111111110001 : data = 16'b1100010111011110;
            15'b000111111110010 : data = 16'b1100010111001101;
            15'b000111111110011 : data = 16'b1100010110111011;
            15'b000111111110100 : data = 16'b1100010110101010;
            15'b000111111110101 : data = 16'b1100010110011001;
            15'b000111111110110 : data = 16'b1100010110001000;
            15'b000111111110111 : data = 16'b1100010101110110;
            15'b000111111111000 : data = 16'b1100010101100101;
            15'b000111111111001 : data = 16'b1100010101010100;
            15'b000111111111010 : data = 16'b1100010101000010;
            15'b000111111111011 : data = 16'b1100010100110001;
            15'b000111111111100 : data = 16'b1100010100100000;
            15'b000111111111101 : data = 16'b1100010100001110;
            15'b000111111111110 : data = 16'b1100010011111101;
            15'b000111111111111 : data = 16'b1100010011101100;
            15'b001000000000000 : data = 16'b1100010011011010;
            15'b001000000000001 : data = 16'b1100010011001001;
            15'b001000000000010 : data = 16'b1100010010111000;
            15'b001000000000011 : data = 16'b1100010010100110;
            15'b001000000000100 : data = 16'b1100010010010101;
            15'b001000000000101 : data = 16'b1100010010000100;
            15'b001000000000110 : data = 16'b1100010001110010;
            15'b001000000000111 : data = 16'b1100010001100001;
            15'b001000000001000 : data = 16'b1100010001001111;
            15'b001000000001001 : data = 16'b1100010000111110;
            15'b001000000001010 : data = 16'b1100010000101101;
            15'b001000000001011 : data = 16'b1100010000011011;
            15'b001000000001100 : data = 16'b1100010000001010;
            15'b001000000001101 : data = 16'b1100001111111000;
            15'b001000000001110 : data = 16'b1100001111100111;
            15'b001000000001111 : data = 16'b1100001111010101;
            15'b001000000010000 : data = 16'b1100001111000100;
            15'b001000000010001 : data = 16'b1100001110110010;
            15'b001000000010010 : data = 16'b1100001110100001;
            15'b001000000010011 : data = 16'b1100001110001111;
            15'b001000000010100 : data = 16'b1100001101111110;
            15'b001000000010101 : data = 16'b1100001101101100;
            15'b001000000010110 : data = 16'b1100001101011011;
            15'b001000000010111 : data = 16'b1100001101001001;
            15'b001000000011000 : data = 16'b1100001100111000;
            15'b001000000011001 : data = 16'b1100001100100110;
            15'b001000000011010 : data = 16'b1100001100010101;
            15'b001000000011011 : data = 16'b1100001100000011;
            15'b001000000011100 : data = 16'b1100001011110010;
            15'b001000000011101 : data = 16'b1100001011100000;
            15'b001000000011110 : data = 16'b1100001011001111;
            15'b001000000011111 : data = 16'b1100001010111101;
            15'b001000000100000 : data = 16'b1100001010101100;
            15'b001000000100001 : data = 16'b1100001010011010;
            15'b001000000100010 : data = 16'b1100001010001000;
            15'b001000000100011 : data = 16'b1100001001110111;
            15'b001000000100100 : data = 16'b1100001001100101;
            15'b001000000100101 : data = 16'b1100001001010100;
            15'b001000000100110 : data = 16'b1100001001000010;
            15'b001000000100111 : data = 16'b1100001000110000;
            15'b001000000101000 : data = 16'b1100001000011111;
            15'b001000000101001 : data = 16'b1100001000001101;
            15'b001000000101010 : data = 16'b1100000111111011;
            15'b001000000101011 : data = 16'b1100000111101010;
            15'b001000000101100 : data = 16'b1100000111011000;
            15'b001000000101101 : data = 16'b1100000111000110;
            15'b001000000101110 : data = 16'b1100000110110101;
            15'b001000000101111 : data = 16'b1100000110100011;
            15'b001000000110000 : data = 16'b1100000110010001;
            15'b001000000110001 : data = 16'b1100000110000000;
            15'b001000000110010 : data = 16'b1100000101101110;
            15'b001000000110011 : data = 16'b1100000101011100;
            15'b001000000110100 : data = 16'b1100000101001011;
            15'b001000000110101 : data = 16'b1100000100111001;
            15'b001000000110110 : data = 16'b1100000100100111;
            15'b001000000110111 : data = 16'b1100000100010110;
            15'b001000000111000 : data = 16'b1100000100000100;
            15'b001000000111001 : data = 16'b1100000011110010;
            15'b001000000111010 : data = 16'b1100000011100000;
            15'b001000000111011 : data = 16'b1100000011001111;
            15'b001000000111100 : data = 16'b1100000010111101;
            15'b001000000111101 : data = 16'b1100000010101011;
            15'b001000000111110 : data = 16'b1100000010011001;
            15'b001000000111111 : data = 16'b1100000010001000;
            15'b001000001000000 : data = 16'b1100000001110110;
            15'b001000001000001 : data = 16'b1100000001100100;
            15'b001000001000010 : data = 16'b1100000001010010;
            15'b001000001000011 : data = 16'b1100000001000000;
            15'b001000001000100 : data = 16'b1100000000101111;
            15'b001000001000101 : data = 16'b1100000000011101;
            15'b001000001000110 : data = 16'b1100000000001011;
            15'b001000001000111 : data = 16'b1011111111111001;
            15'b001000001001000 : data = 16'b1011111111100111;
            15'b001000001001001 : data = 16'b1011111111010101;
            15'b001000001001010 : data = 16'b1011111111000100;
            15'b001000001001011 : data = 16'b1011111110110010;
            15'b001000001001100 : data = 16'b1011111110100000;
            15'b001000001001101 : data = 16'b1011111110001110;
            15'b001000001001110 : data = 16'b1011111101111100;
            15'b001000001001111 : data = 16'b1011111101101010;
            15'b001000001010000 : data = 16'b1011111101011000;
            15'b001000001010001 : data = 16'b1011111101000110;
            15'b001000001010010 : data = 16'b1011111100110101;
            15'b001000001010011 : data = 16'b1011111100100011;
            15'b001000001010100 : data = 16'b1011111100010001;
            15'b001000001010101 : data = 16'b1011111011111111;
            15'b001000001010110 : data = 16'b1011111011101101;
            15'b001000001010111 : data = 16'b1011111011011011;
            15'b001000001011000 : data = 16'b1011111011001001;
            15'b001000001011001 : data = 16'b1011111010110111;
            15'b001000001011010 : data = 16'b1011111010100101;
            15'b001000001011011 : data = 16'b1011111010010011;
            15'b001000001011100 : data = 16'b1011111010000001;
            15'b001000001011101 : data = 16'b1011111001101111;
            15'b001000001011110 : data = 16'b1011111001011101;
            15'b001000001011111 : data = 16'b1011111001001011;
            15'b001000001100000 : data = 16'b1011111000111001;
            15'b001000001100001 : data = 16'b1011111000100111;
            15'b001000001100010 : data = 16'b1011111000010101;
            15'b001000001100011 : data = 16'b1011111000000011;
            15'b001000001100100 : data = 16'b1011110111110001;
            15'b001000001100101 : data = 16'b1011110111011111;
            15'b001000001100110 : data = 16'b1011110111001101;
            15'b001000001100111 : data = 16'b1011110110111011;
            15'b001000001101000 : data = 16'b1011110110101001;
            15'b001000001101001 : data = 16'b1011110110010111;
            15'b001000001101010 : data = 16'b1011110110000101;
            15'b001000001101011 : data = 16'b1011110101110011;
            15'b001000001101100 : data = 16'b1011110101100001;
            15'b001000001101101 : data = 16'b1011110101001111;
            15'b001000001101110 : data = 16'b1011110100111101;
            15'b001000001101111 : data = 16'b1011110100101011;
            15'b001000001110000 : data = 16'b1011110100011001;
            15'b001000001110001 : data = 16'b1011110100000110;
            15'b001000001110010 : data = 16'b1011110011110100;
            15'b001000001110011 : data = 16'b1011110011100010;
            15'b001000001110100 : data = 16'b1011110011010000;
            15'b001000001110101 : data = 16'b1011110010111110;
            15'b001000001110110 : data = 16'b1011110010101100;
            15'b001000001110111 : data = 16'b1011110010011010;
            15'b001000001111000 : data = 16'b1011110010001000;
            15'b001000001111001 : data = 16'b1011110001110110;
            15'b001000001111010 : data = 16'b1011110001100011;
            15'b001000001111011 : data = 16'b1011110001010001;
            15'b001000001111100 : data = 16'b1011110000111111;
            15'b001000001111101 : data = 16'b1011110000101101;
            15'b001000001111110 : data = 16'b1011110000011011;
            15'b001000001111111 : data = 16'b1011110000001001;
            15'b001000010000000 : data = 16'b1011101111110110;
            15'b001000010000001 : data = 16'b1011101111100100;
            15'b001000010000010 : data = 16'b1011101111010010;
            15'b001000010000011 : data = 16'b1011101111000000;
            15'b001000010000100 : data = 16'b1011101110101110;
            15'b001000010000101 : data = 16'b1011101110011011;
            15'b001000010000110 : data = 16'b1011101110001001;
            15'b001000010000111 : data = 16'b1011101101110111;
            15'b001000010001000 : data = 16'b1011101101100101;
            15'b001000010001001 : data = 16'b1011101101010010;
            15'b001000010001010 : data = 16'b1011101101000000;
            15'b001000010001011 : data = 16'b1011101100101110;
            15'b001000010001100 : data = 16'b1011101100011100;
            15'b001000010001101 : data = 16'b1011101100001001;
            15'b001000010001110 : data = 16'b1011101011110111;
            15'b001000010001111 : data = 16'b1011101011100101;
            15'b001000010010000 : data = 16'b1011101011010011;
            15'b001000010010001 : data = 16'b1011101011000000;
            15'b001000010010010 : data = 16'b1011101010101110;
            15'b001000010010011 : data = 16'b1011101010011100;
            15'b001000010010100 : data = 16'b1011101010001001;
            15'b001000010010101 : data = 16'b1011101001110111;
            15'b001000010010110 : data = 16'b1011101001100101;
            15'b001000010010111 : data = 16'b1011101001010010;
            15'b001000010011000 : data = 16'b1011101001000000;
            15'b001000010011001 : data = 16'b1011101000101110;
            15'b001000010011010 : data = 16'b1011101000011011;
            15'b001000010011011 : data = 16'b1011101000001001;
            15'b001000010011100 : data = 16'b1011100111110111;
            15'b001000010011101 : data = 16'b1011100111100100;
            15'b001000010011110 : data = 16'b1011100111010010;
            15'b001000010011111 : data = 16'b1011100111000000;
            15'b001000010100000 : data = 16'b1011100110101101;
            15'b001000010100001 : data = 16'b1011100110011011;
            15'b001000010100010 : data = 16'b1011100110001000;
            15'b001000010100011 : data = 16'b1011100101110110;
            15'b001000010100100 : data = 16'b1011100101100100;
            15'b001000010100101 : data = 16'b1011100101010001;
            15'b001000010100110 : data = 16'b1011100100111111;
            15'b001000010100111 : data = 16'b1011100100101100;
            15'b001000010101000 : data = 16'b1011100100011010;
            15'b001000010101001 : data = 16'b1011100100001000;
            15'b001000010101010 : data = 16'b1011100011110101;
            15'b001000010101011 : data = 16'b1011100011100011;
            15'b001000010101100 : data = 16'b1011100011010000;
            15'b001000010101101 : data = 16'b1011100010111110;
            15'b001000010101110 : data = 16'b1011100010101011;
            15'b001000010101111 : data = 16'b1011100010011001;
            15'b001000010110000 : data = 16'b1011100010000110;
            15'b001000010110001 : data = 16'b1011100001110100;
            15'b001000010110010 : data = 16'b1011100001100001;
            15'b001000010110011 : data = 16'b1011100001001111;
            15'b001000010110100 : data = 16'b1011100000111100;
            15'b001000010110101 : data = 16'b1011100000101010;
            15'b001000010110110 : data = 16'b1011100000010111;
            15'b001000010110111 : data = 16'b1011100000000101;
            15'b001000010111000 : data = 16'b1011011111110010;
            15'b001000010111001 : data = 16'b1011011111100000;
            15'b001000010111010 : data = 16'b1011011111001101;
            15'b001000010111011 : data = 16'b1011011110111011;
            15'b001000010111100 : data = 16'b1011011110101000;
            15'b001000010111101 : data = 16'b1011011110010110;
            15'b001000010111110 : data = 16'b1011011110000011;
            15'b001000010111111 : data = 16'b1011011101110001;
            15'b001000011000000 : data = 16'b1011011101011110;
            15'b001000011000001 : data = 16'b1011011101001100;
            15'b001000011000010 : data = 16'b1011011100111001;
            15'b001000011000011 : data = 16'b1011011100100110;
            15'b001000011000100 : data = 16'b1011011100010100;
            15'b001000011000101 : data = 16'b1011011100000001;
            15'b001000011000110 : data = 16'b1011011011101111;
            15'b001000011000111 : data = 16'b1011011011011100;
            15'b001000011001000 : data = 16'b1011011011001001;
            15'b001000011001001 : data = 16'b1011011010110111;
            15'b001000011001010 : data = 16'b1011011010100100;
            15'b001000011001011 : data = 16'b1011011010010010;
            15'b001000011001100 : data = 16'b1011011001111111;
            15'b001000011001101 : data = 16'b1011011001101100;
            15'b001000011001110 : data = 16'b1011011001011010;
            15'b001000011001111 : data = 16'b1011011001000111;
            15'b001000011010000 : data = 16'b1011011000110100;
            15'b001000011010001 : data = 16'b1011011000100010;
            15'b001000011010010 : data = 16'b1011011000001111;
            15'b001000011010011 : data = 16'b1011010111111100;
            15'b001000011010100 : data = 16'b1011010111101010;
            15'b001000011010101 : data = 16'b1011010111010111;
            15'b001000011010110 : data = 16'b1011010111000100;
            15'b001000011010111 : data = 16'b1011010110110010;
            15'b001000011011000 : data = 16'b1011010110011111;
            15'b001000011011001 : data = 16'b1011010110001100;
            15'b001000011011010 : data = 16'b1011010101111010;
            15'b001000011011011 : data = 16'b1011010101100111;
            15'b001000011011100 : data = 16'b1011010101010100;
            15'b001000011011101 : data = 16'b1011010101000010;
            15'b001000011011110 : data = 16'b1011010100101111;
            15'b001000011011111 : data = 16'b1011010100011100;
            15'b001000011100000 : data = 16'b1011010100001001;
            15'b001000011100001 : data = 16'b1011010011110111;
            15'b001000011100010 : data = 16'b1011010011100100;
            15'b001000011100011 : data = 16'b1011010011010001;
            15'b001000011100100 : data = 16'b1011010010111110;
            15'b001000011100101 : data = 16'b1011010010101100;
            15'b001000011100110 : data = 16'b1011010010011001;
            15'b001000011100111 : data = 16'b1011010010000110;
            15'b001000011101000 : data = 16'b1011010001110011;
            15'b001000011101001 : data = 16'b1011010001100000;
            15'b001000011101010 : data = 16'b1011010001001110;
            15'b001000011101011 : data = 16'b1011010000111011;
            15'b001000011101100 : data = 16'b1011010000101000;
            15'b001000011101101 : data = 16'b1011010000010101;
            15'b001000011101110 : data = 16'b1011010000000010;
            15'b001000011101111 : data = 16'b1011001111110000;
            15'b001000011110000 : data = 16'b1011001111011101;
            15'b001000011110001 : data = 16'b1011001111001010;
            15'b001000011110010 : data = 16'b1011001110110111;
            15'b001000011110011 : data = 16'b1011001110100100;
            15'b001000011110100 : data = 16'b1011001110010010;
            15'b001000011110101 : data = 16'b1011001101111111;
            15'b001000011110110 : data = 16'b1011001101101100;
            15'b001000011110111 : data = 16'b1011001101011001;
            15'b001000011111000 : data = 16'b1011001101000110;
            15'b001000011111001 : data = 16'b1011001100110011;
            15'b001000011111010 : data = 16'b1011001100100000;
            15'b001000011111011 : data = 16'b1011001100001110;
            15'b001000011111100 : data = 16'b1011001011111011;
            15'b001000011111101 : data = 16'b1011001011101000;
            15'b001000011111110 : data = 16'b1011001011010101;
            15'b001000011111111 : data = 16'b1011001011000010;
            15'b001000100000000 : data = 16'b1011001010101111;
            15'b001000100000001 : data = 16'b1011001010011100;
            15'b001000100000010 : data = 16'b1011001010001001;
            15'b001000100000011 : data = 16'b1011001001110110;
            15'b001000100000100 : data = 16'b1011001001100011;
            15'b001000100000101 : data = 16'b1011001001010000;
            15'b001000100000110 : data = 16'b1011001000111110;
            15'b001000100000111 : data = 16'b1011001000101011;
            15'b001000100001000 : data = 16'b1011001000011000;
            15'b001000100001001 : data = 16'b1011001000000101;
            15'b001000100001010 : data = 16'b1011000111110010;
            15'b001000100001011 : data = 16'b1011000111011111;
            15'b001000100001100 : data = 16'b1011000111001100;
            15'b001000100001101 : data = 16'b1011000110111001;
            15'b001000100001110 : data = 16'b1011000110100110;
            15'b001000100001111 : data = 16'b1011000110010011;
            15'b001000100010000 : data = 16'b1011000110000000;
            15'b001000100010001 : data = 16'b1011000101101101;
            15'b001000100010010 : data = 16'b1011000101011010;
            15'b001000100010011 : data = 16'b1011000101000111;
            15'b001000100010100 : data = 16'b1011000100110100;
            15'b001000100010101 : data = 16'b1011000100100001;
            15'b001000100010110 : data = 16'b1011000100001110;
            15'b001000100010111 : data = 16'b1011000011111011;
            15'b001000100011000 : data = 16'b1011000011101000;
            15'b001000100011001 : data = 16'b1011000011010101;
            15'b001000100011010 : data = 16'b1011000011000010;
            15'b001000100011011 : data = 16'b1011000010101111;
            15'b001000100011100 : data = 16'b1011000010011100;
            15'b001000100011101 : data = 16'b1011000010001001;
            15'b001000100011110 : data = 16'b1011000001110110;
            15'b001000100011111 : data = 16'b1011000001100011;
            15'b001000100100000 : data = 16'b1011000001010000;
            15'b001000100100001 : data = 16'b1011000000111100;
            15'b001000100100010 : data = 16'b1011000000101001;
            15'b001000100100011 : data = 16'b1011000000010110;
            15'b001000100100100 : data = 16'b1011000000000011;
            15'b001000100100101 : data = 16'b1010111111110000;
            15'b001000100100110 : data = 16'b1010111111011101;
            15'b001000100100111 : data = 16'b1010111111001010;
            15'b001000100101000 : data = 16'b1010111110110111;
            15'b001000100101001 : data = 16'b1010111110100100;
            15'b001000100101010 : data = 16'b1010111110010001;
            15'b001000100101011 : data = 16'b1010111101111101;
            15'b001000100101100 : data = 16'b1010111101101010;
            15'b001000100101101 : data = 16'b1010111101010111;
            15'b001000100101110 : data = 16'b1010111101000100;
            15'b001000100101111 : data = 16'b1010111100110001;
            15'b001000100110000 : data = 16'b1010111100011110;
            15'b001000100110001 : data = 16'b1010111100001011;
            15'b001000100110010 : data = 16'b1010111011111000;
            15'b001000100110011 : data = 16'b1010111011100100;
            15'b001000100110100 : data = 16'b1010111011010001;
            15'b001000100110101 : data = 16'b1010111010111110;
            15'b001000100110110 : data = 16'b1010111010101011;
            15'b001000100110111 : data = 16'b1010111010011000;
            15'b001000100111000 : data = 16'b1010111010000101;
            15'b001000100111001 : data = 16'b1010111001110001;
            15'b001000100111010 : data = 16'b1010111001011110;
            15'b001000100111011 : data = 16'b1010111001001011;
            15'b001000100111100 : data = 16'b1010111000111000;
            15'b001000100111101 : data = 16'b1010111000100101;
            15'b001000100111110 : data = 16'b1010111000010001;
            15'b001000100111111 : data = 16'b1010110111111110;
            15'b001000101000000 : data = 16'b1010110111101011;
            15'b001000101000001 : data = 16'b1010110111011000;
            15'b001000101000010 : data = 16'b1010110111000101;
            15'b001000101000011 : data = 16'b1010110110110001;
            15'b001000101000100 : data = 16'b1010110110011110;
            15'b001000101000101 : data = 16'b1010110110001011;
            15'b001000101000110 : data = 16'b1010110101111000;
            15'b001000101000111 : data = 16'b1010110101100100;
            15'b001000101001000 : data = 16'b1010110101010001;
            15'b001000101001001 : data = 16'b1010110100111110;
            15'b001000101001010 : data = 16'b1010110100101011;
            15'b001000101001011 : data = 16'b1010110100010111;
            15'b001000101001100 : data = 16'b1010110100000100;
            15'b001000101001101 : data = 16'b1010110011110001;
            15'b001000101001110 : data = 16'b1010110011011101;
            15'b001000101001111 : data = 16'b1010110011001010;
            15'b001000101010000 : data = 16'b1010110010110111;
            15'b001000101010001 : data = 16'b1010110010100100;
            15'b001000101010010 : data = 16'b1010110010010000;
            15'b001000101010011 : data = 16'b1010110001111101;
            15'b001000101010100 : data = 16'b1010110001101010;
            15'b001000101010101 : data = 16'b1010110001010110;
            15'b001000101010110 : data = 16'b1010110001000011;
            15'b001000101010111 : data = 16'b1010110000110000;
            15'b001000101011000 : data = 16'b1010110000011100;
            15'b001000101011001 : data = 16'b1010110000001001;
            15'b001000101011010 : data = 16'b1010101111110110;
            15'b001000101011011 : data = 16'b1010101111100010;
            15'b001000101011100 : data = 16'b1010101111001111;
            15'b001000101011101 : data = 16'b1010101110111100;
            15'b001000101011110 : data = 16'b1010101110101000;
            15'b001000101011111 : data = 16'b1010101110010101;
            15'b001000101100000 : data = 16'b1010101110000010;
            15'b001000101100001 : data = 16'b1010101101101110;
            15'b001000101100010 : data = 16'b1010101101011011;
            15'b001000101100011 : data = 16'b1010101101001000;
            15'b001000101100100 : data = 16'b1010101100110100;
            15'b001000101100101 : data = 16'b1010101100100001;
            15'b001000101100110 : data = 16'b1010101100001101;
            15'b001000101100111 : data = 16'b1010101011111010;
            15'b001000101101000 : data = 16'b1010101011100111;
            15'b001000101101001 : data = 16'b1010101011010011;
            15'b001000101101010 : data = 16'b1010101011000000;
            15'b001000101101011 : data = 16'b1010101010101100;
            15'b001000101101100 : data = 16'b1010101010011001;
            15'b001000101101101 : data = 16'b1010101010000110;
            15'b001000101101110 : data = 16'b1010101001110010;
            15'b001000101101111 : data = 16'b1010101001011111;
            15'b001000101110000 : data = 16'b1010101001001011;
            15'b001000101110001 : data = 16'b1010101000111000;
            15'b001000101110010 : data = 16'b1010101000100100;
            15'b001000101110011 : data = 16'b1010101000010001;
            15'b001000101110100 : data = 16'b1010100111111110;
            15'b001000101110101 : data = 16'b1010100111101010;
            15'b001000101110110 : data = 16'b1010100111010111;
            15'b001000101110111 : data = 16'b1010100111000011;
            15'b001000101111000 : data = 16'b1010100110110000;
            15'b001000101111001 : data = 16'b1010100110011100;
            15'b001000101111010 : data = 16'b1010100110001001;
            15'b001000101111011 : data = 16'b1010100101110101;
            15'b001000101111100 : data = 16'b1010100101100010;
            15'b001000101111101 : data = 16'b1010100101001110;
            15'b001000101111110 : data = 16'b1010100100111011;
            15'b001000101111111 : data = 16'b1010100100100111;
            15'b001000110000000 : data = 16'b1010100100010100;
            15'b001000110000001 : data = 16'b1010100100000000;
            15'b001000110000010 : data = 16'b1010100011101101;
            15'b001000110000011 : data = 16'b1010100011011001;
            15'b001000110000100 : data = 16'b1010100011000110;
            15'b001000110000101 : data = 16'b1010100010110010;
            15'b001000110000110 : data = 16'b1010100010011111;
            15'b001000110000111 : data = 16'b1010100010001011;
            15'b001000110001000 : data = 16'b1010100001111000;
            15'b001000110001001 : data = 16'b1010100001100100;
            15'b001000110001010 : data = 16'b1010100001010001;
            15'b001000110001011 : data = 16'b1010100000111101;
            15'b001000110001100 : data = 16'b1010100000101010;
            15'b001000110001101 : data = 16'b1010100000010110;
            15'b001000110001110 : data = 16'b1010100000000010;
            15'b001000110001111 : data = 16'b1010011111101111;
            15'b001000110010000 : data = 16'b1010011111011011;
            15'b001000110010001 : data = 16'b1010011111001000;
            15'b001000110010010 : data = 16'b1010011110110100;
            15'b001000110010011 : data = 16'b1010011110100001;
            15'b001000110010100 : data = 16'b1010011110001101;
            15'b001000110010101 : data = 16'b1010011101111001;
            15'b001000110010110 : data = 16'b1010011101100110;
            15'b001000110010111 : data = 16'b1010011101010010;
            15'b001000110011000 : data = 16'b1010011100111111;
            15'b001000110011001 : data = 16'b1010011100101011;
            15'b001000110011010 : data = 16'b1010011100011000;
            15'b001000110011011 : data = 16'b1010011100000100;
            15'b001000110011100 : data = 16'b1010011011110000;
            15'b001000110011101 : data = 16'b1010011011011101;
            15'b001000110011110 : data = 16'b1010011011001001;
            15'b001000110011111 : data = 16'b1010011010110101;
            15'b001000110100000 : data = 16'b1010011010100010;
            15'b001000110100001 : data = 16'b1010011010001110;
            15'b001000110100010 : data = 16'b1010011001111011;
            15'b001000110100011 : data = 16'b1010011001100111;
            15'b001000110100100 : data = 16'b1010011001010011;
            15'b001000110100101 : data = 16'b1010011001000000;
            15'b001000110100110 : data = 16'b1010011000101100;
            15'b001000110100111 : data = 16'b1010011000011000;
            15'b001000110101000 : data = 16'b1010011000000101;
            15'b001000110101001 : data = 16'b1010010111110001;
            15'b001000110101010 : data = 16'b1010010111011101;
            15'b001000110101011 : data = 16'b1010010111001010;
            15'b001000110101100 : data = 16'b1010010110110110;
            15'b001000110101101 : data = 16'b1010010110100010;
            15'b001000110101110 : data = 16'b1010010110001111;
            15'b001000110101111 : data = 16'b1010010101111011;
            15'b001000110110000 : data = 16'b1010010101100111;
            15'b001000110110001 : data = 16'b1010010101010100;
            15'b001000110110010 : data = 16'b1010010101000000;
            15'b001000110110011 : data = 16'b1010010100101100;
            15'b001000110110100 : data = 16'b1010010100011000;
            15'b001000110110101 : data = 16'b1010010100000101;
            15'b001000110110110 : data = 16'b1010010011110001;
            15'b001000110110111 : data = 16'b1010010011011101;
            15'b001000110111000 : data = 16'b1010010011001010;
            15'b001000110111001 : data = 16'b1010010010110110;
            15'b001000110111010 : data = 16'b1010010010100010;
            15'b001000110111011 : data = 16'b1010010010001110;
            15'b001000110111100 : data = 16'b1010010001111011;
            15'b001000110111101 : data = 16'b1010010001100111;
            15'b001000110111110 : data = 16'b1010010001010011;
            15'b001000110111111 : data = 16'b1010010001000000;
            15'b001000111000000 : data = 16'b1010010000101100;
            15'b001000111000001 : data = 16'b1010010000011000;
            15'b001000111000010 : data = 16'b1010010000000100;
            15'b001000111000011 : data = 16'b1010001111110000;
            15'b001000111000100 : data = 16'b1010001111011101;
            15'b001000111000101 : data = 16'b1010001111001001;
            15'b001000111000110 : data = 16'b1010001110110101;
            15'b001000111000111 : data = 16'b1010001110100001;
            15'b001000111001000 : data = 16'b1010001110001110;
            15'b001000111001001 : data = 16'b1010001101111010;
            15'b001000111001010 : data = 16'b1010001101100110;
            15'b001000111001011 : data = 16'b1010001101010010;
            15'b001000111001100 : data = 16'b1010001100111111;
            15'b001000111001101 : data = 16'b1010001100101011;
            15'b001000111001110 : data = 16'b1010001100010111;
            15'b001000111001111 : data = 16'b1010001100000011;
            15'b001000111010000 : data = 16'b1010001011101111;
            15'b001000111010001 : data = 16'b1010001011011100;
            15'b001000111010010 : data = 16'b1010001011001000;
            15'b001000111010011 : data = 16'b1010001010110100;
            15'b001000111010100 : data = 16'b1010001010100000;
            15'b001000111010101 : data = 16'b1010001010001100;
            15'b001000111010110 : data = 16'b1010001001111000;
            15'b001000111010111 : data = 16'b1010001001100101;
            15'b001000111011000 : data = 16'b1010001001010001;
            15'b001000111011001 : data = 16'b1010001000111101;
            15'b001000111011010 : data = 16'b1010001000101001;
            15'b001000111011011 : data = 16'b1010001000010101;
            15'b001000111011100 : data = 16'b1010001000000001;
            15'b001000111011101 : data = 16'b1010000111101110;
            15'b001000111011110 : data = 16'b1010000111011010;
            15'b001000111011111 : data = 16'b1010000111000110;
            15'b001000111100000 : data = 16'b1010000110110010;
            15'b001000111100001 : data = 16'b1010000110011110;
            15'b001000111100010 : data = 16'b1010000110001010;
            15'b001000111100011 : data = 16'b1010000101110110;
            15'b001000111100100 : data = 16'b1010000101100010;
            15'b001000111100101 : data = 16'b1010000101001111;
            15'b001000111100110 : data = 16'b1010000100111011;
            15'b001000111100111 : data = 16'b1010000100100111;
            15'b001000111101000 : data = 16'b1010000100010011;
            15'b001000111101001 : data = 16'b1010000011111111;
            15'b001000111101010 : data = 16'b1010000011101011;
            15'b001000111101011 : data = 16'b1010000011010111;
            15'b001000111101100 : data = 16'b1010000011000011;
            15'b001000111101101 : data = 16'b1010000010101111;
            15'b001000111101110 : data = 16'b1010000010011100;
            15'b001000111101111 : data = 16'b1010000010001000;
            15'b001000111110000 : data = 16'b1010000001110100;
            15'b001000111110001 : data = 16'b1010000001100000;
            15'b001000111110010 : data = 16'b1010000001001100;
            15'b001000111110011 : data = 16'b1010000000111000;
            15'b001000111110100 : data = 16'b1010000000100100;
            15'b001000111110101 : data = 16'b1010000000010000;
            15'b001000111110110 : data = 16'b1001111111111100;
            15'b001000111110111 : data = 16'b1001111111101000;
            15'b001000111111000 : data = 16'b1001111111010100;
            15'b001000111111001 : data = 16'b1001111111000000;
            15'b001000111111010 : data = 16'b1001111110101100;
            15'b001000111111011 : data = 16'b1001111110011000;
            15'b001000111111100 : data = 16'b1001111110000101;
            15'b001000111111101 : data = 16'b1001111101110001;
            15'b001000111111110 : data = 16'b1001111101011101;
            15'b001000111111111 : data = 16'b1001111101001001;
            15'b001001000000000 : data = 16'b1001111100110101;
            15'b001001000000001 : data = 16'b1001111100100001;
            15'b001001000000010 : data = 16'b1001111100001101;
            15'b001001000000011 : data = 16'b1001111011111001;
            15'b001001000000100 : data = 16'b1001111011100101;
            15'b001001000000101 : data = 16'b1001111011010001;
            15'b001001000000110 : data = 16'b1001111010111101;
            15'b001001000000111 : data = 16'b1001111010101001;
            15'b001001000001000 : data = 16'b1001111010010101;
            15'b001001000001001 : data = 16'b1001111010000001;
            15'b001001000001010 : data = 16'b1001111001101101;
            15'b001001000001011 : data = 16'b1001111001011001;
            15'b001001000001100 : data = 16'b1001111001000101;
            15'b001001000001101 : data = 16'b1001111000110001;
            15'b001001000001110 : data = 16'b1001111000011101;
            15'b001001000001111 : data = 16'b1001111000001001;
            15'b001001000010000 : data = 16'b1001110111110101;
            15'b001001000010001 : data = 16'b1001110111100001;
            15'b001001000010010 : data = 16'b1001110111001101;
            15'b001001000010011 : data = 16'b1001110110111001;
            15'b001001000010100 : data = 16'b1001110110100101;
            15'b001001000010101 : data = 16'b1001110110010001;
            15'b001001000010110 : data = 16'b1001110101111101;
            15'b001001000010111 : data = 16'b1001110101101001;
            15'b001001000011000 : data = 16'b1001110101010101;
            15'b001001000011001 : data = 16'b1001110101000001;
            15'b001001000011010 : data = 16'b1001110100101101;
            15'b001001000011011 : data = 16'b1001110100011000;
            15'b001001000011100 : data = 16'b1001110100000100;
            15'b001001000011101 : data = 16'b1001110011110000;
            15'b001001000011110 : data = 16'b1001110011011100;
            15'b001001000011111 : data = 16'b1001110011001000;
            15'b001001000100000 : data = 16'b1001110010110100;
            15'b001001000100001 : data = 16'b1001110010100000;
            15'b001001000100010 : data = 16'b1001110010001100;
            15'b001001000100011 : data = 16'b1001110001111000;
            15'b001001000100100 : data = 16'b1001110001100100;
            15'b001001000100101 : data = 16'b1001110001010000;
            15'b001001000100110 : data = 16'b1001110000111100;
            15'b001001000100111 : data = 16'b1001110000101000;
            15'b001001000101000 : data = 16'b1001110000010100;
            15'b001001000101001 : data = 16'b1001101111111111;
            15'b001001000101010 : data = 16'b1001101111101011;
            15'b001001000101011 : data = 16'b1001101111010111;
            15'b001001000101100 : data = 16'b1001101111000011;
            15'b001001000101101 : data = 16'b1001101110101111;
            15'b001001000101110 : data = 16'b1001101110011011;
            15'b001001000101111 : data = 16'b1001101110000111;
            15'b001001000110000 : data = 16'b1001101101110011;
            15'b001001000110001 : data = 16'b1001101101011111;
            15'b001001000110010 : data = 16'b1001101101001011;
            15'b001001000110011 : data = 16'b1001101100110110;
            15'b001001000110100 : data = 16'b1001101100100010;
            15'b001001000110101 : data = 16'b1001101100001110;
            15'b001001000110110 : data = 16'b1001101011111010;
            15'b001001000110111 : data = 16'b1001101011100110;
            15'b001001000111000 : data = 16'b1001101011010010;
            15'b001001000111001 : data = 16'b1001101010111110;
            15'b001001000111010 : data = 16'b1001101010101010;
            15'b001001000111011 : data = 16'b1001101010010101;
            15'b001001000111100 : data = 16'b1001101010000001;
            15'b001001000111101 : data = 16'b1001101001101101;
            15'b001001000111110 : data = 16'b1001101001011001;
            15'b001001000111111 : data = 16'b1001101001000101;
            15'b001001001000000 : data = 16'b1001101000110001;
            15'b001001001000001 : data = 16'b1001101000011101;
            15'b001001001000010 : data = 16'b1001101000001000;
            15'b001001001000011 : data = 16'b1001100111110100;
            15'b001001001000100 : data = 16'b1001100111100000;
            15'b001001001000101 : data = 16'b1001100111001100;
            15'b001001001000110 : data = 16'b1001100110111000;
            15'b001001001000111 : data = 16'b1001100110100100;
            15'b001001001001000 : data = 16'b1001100110001111;
            15'b001001001001001 : data = 16'b1001100101111011;
            15'b001001001001010 : data = 16'b1001100101100111;
            15'b001001001001011 : data = 16'b1001100101010011;
            15'b001001001001100 : data = 16'b1001100100111111;
            15'b001001001001101 : data = 16'b1001100100101010;
            15'b001001001001110 : data = 16'b1001100100010110;
            15'b001001001001111 : data = 16'b1001100100000010;
            15'b001001001010000 : data = 16'b1001100011101110;
            15'b001001001010001 : data = 16'b1001100011011010;
            15'b001001001010010 : data = 16'b1001100011000110;
            15'b001001001010011 : data = 16'b1001100010110001;
            15'b001001001010100 : data = 16'b1001100010011101;
            15'b001001001010101 : data = 16'b1001100010001001;
            15'b001001001010110 : data = 16'b1001100001110101;
            15'b001001001010111 : data = 16'b1001100001100001;
            15'b001001001011000 : data = 16'b1001100001001100;
            15'b001001001011001 : data = 16'b1001100000111000;
            15'b001001001011010 : data = 16'b1001100000100100;
            15'b001001001011011 : data = 16'b1001100000010000;
            15'b001001001011100 : data = 16'b1001011111111011;
            15'b001001001011101 : data = 16'b1001011111100111;
            15'b001001001011110 : data = 16'b1001011111010011;
            15'b001001001011111 : data = 16'b1001011110111111;
            15'b001001001100000 : data = 16'b1001011110101011;
            15'b001001001100001 : data = 16'b1001011110010110;
            15'b001001001100010 : data = 16'b1001011110000010;
            15'b001001001100011 : data = 16'b1001011101101110;
            15'b001001001100100 : data = 16'b1001011101011010;
            15'b001001001100101 : data = 16'b1001011101000101;
            15'b001001001100110 : data = 16'b1001011100110001;
            15'b001001001100111 : data = 16'b1001011100011101;
            15'b001001001101000 : data = 16'b1001011100001001;
            15'b001001001101001 : data = 16'b1001011011110100;
            15'b001001001101010 : data = 16'b1001011011100000;
            15'b001001001101011 : data = 16'b1001011011001100;
            15'b001001001101100 : data = 16'b1001011010111000;
            15'b001001001101101 : data = 16'b1001011010100011;
            15'b001001001101110 : data = 16'b1001011010001111;
            15'b001001001101111 : data = 16'b1001011001111011;
            15'b001001001110000 : data = 16'b1001011001100110;
            15'b001001001110001 : data = 16'b1001011001010010;
            15'b001001001110010 : data = 16'b1001011000111110;
            15'b001001001110011 : data = 16'b1001011000101010;
            15'b001001001110100 : data = 16'b1001011000010101;
            15'b001001001110101 : data = 16'b1001011000000001;
            15'b001001001110110 : data = 16'b1001010111101101;
            15'b001001001110111 : data = 16'b1001010111011001;
            15'b001001001111000 : data = 16'b1001010111000100;
            15'b001001001111001 : data = 16'b1001010110110000;
            15'b001001001111010 : data = 16'b1001010110011100;
            15'b001001001111011 : data = 16'b1001010110000111;
            15'b001001001111100 : data = 16'b1001010101110011;
            15'b001001001111101 : data = 16'b1001010101011111;
            15'b001001001111110 : data = 16'b1001010101001010;
            15'b001001001111111 : data = 16'b1001010100110110;
            15'b001001010000000 : data = 16'b1001010100100010;
            15'b001001010000001 : data = 16'b1001010100001110;
            15'b001001010000010 : data = 16'b1001010011111001;
            15'b001001010000011 : data = 16'b1001010011100101;
            15'b001001010000100 : data = 16'b1001010011010001;
            15'b001001010000101 : data = 16'b1001010010111100;
            15'b001001010000110 : data = 16'b1001010010101000;
            15'b001001010000111 : data = 16'b1001010010010100;
            15'b001001010001000 : data = 16'b1001010001111111;
            15'b001001010001001 : data = 16'b1001010001101011;
            15'b001001010001010 : data = 16'b1001010001010111;
            15'b001001010001011 : data = 16'b1001010001000010;
            15'b001001010001100 : data = 16'b1001010000101110;
            15'b001001010001101 : data = 16'b1001010000011010;
            15'b001001010001110 : data = 16'b1001010000000101;
            15'b001001010001111 : data = 16'b1001001111110001;
            15'b001001010010000 : data = 16'b1001001111011101;
            15'b001001010010001 : data = 16'b1001001111001000;
            15'b001001010010010 : data = 16'b1001001110110100;
            15'b001001010010011 : data = 16'b1001001110100000;
            15'b001001010010100 : data = 16'b1001001110001011;
            15'b001001010010101 : data = 16'b1001001101110111;
            15'b001001010010110 : data = 16'b1001001101100011;
            15'b001001010010111 : data = 16'b1001001101001110;
            15'b001001010011000 : data = 16'b1001001100111010;
            15'b001001010011001 : data = 16'b1001001100100110;
            15'b001001010011010 : data = 16'b1001001100010001;
            15'b001001010011011 : data = 16'b1001001011111101;
            15'b001001010011100 : data = 16'b1001001011101001;
            15'b001001010011101 : data = 16'b1001001011010100;
            15'b001001010011110 : data = 16'b1001001011000000;
            15'b001001010011111 : data = 16'b1001001010101011;
            15'b001001010100000 : data = 16'b1001001010010111;
            15'b001001010100001 : data = 16'b1001001010000011;
            15'b001001010100010 : data = 16'b1001001001101110;
            15'b001001010100011 : data = 16'b1001001001011010;
            15'b001001010100100 : data = 16'b1001001001000110;
            15'b001001010100101 : data = 16'b1001001000110001;
            15'b001001010100110 : data = 16'b1001001000011101;
            15'b001001010100111 : data = 16'b1001001000001000;
            15'b001001010101000 : data = 16'b1001000111110100;
            15'b001001010101001 : data = 16'b1001000111100000;
            15'b001001010101010 : data = 16'b1001000111001011;
            15'b001001010101011 : data = 16'b1001000110110111;
            15'b001001010101100 : data = 16'b1001000110100010;
            15'b001001010101101 : data = 16'b1001000110001110;
            15'b001001010101110 : data = 16'b1001000101111010;
            15'b001001010101111 : data = 16'b1001000101100101;
            15'b001001010110000 : data = 16'b1001000101010001;
            15'b001001010110001 : data = 16'b1001000100111100;
            15'b001001010110010 : data = 16'b1001000100101000;
            15'b001001010110011 : data = 16'b1001000100010100;
            15'b001001010110100 : data = 16'b1001000011111111;
            15'b001001010110101 : data = 16'b1001000011101011;
            15'b001001010110110 : data = 16'b1001000011010110;
            15'b001001010110111 : data = 16'b1001000011000010;
            15'b001001010111000 : data = 16'b1001000010101110;
            15'b001001010111001 : data = 16'b1001000010011001;
            15'b001001010111010 : data = 16'b1001000010000101;
            15'b001001010111011 : data = 16'b1001000001110000;
            15'b001001010111100 : data = 16'b1001000001011100;
            15'b001001010111101 : data = 16'b1001000001001000;
            15'b001001010111110 : data = 16'b1001000000110011;
            15'b001001010111111 : data = 16'b1001000000011111;
            15'b001001011000000 : data = 16'b1001000000001010;
            15'b001001011000001 : data = 16'b1000111111110110;
            15'b001001011000010 : data = 16'b1000111111100001;
            15'b001001011000011 : data = 16'b1000111111001101;
            15'b001001011000100 : data = 16'b1000111110111001;
            15'b001001011000101 : data = 16'b1000111110100100;
            15'b001001011000110 : data = 16'b1000111110010000;
            15'b001001011000111 : data = 16'b1000111101111011;
            15'b001001011001000 : data = 16'b1000111101100111;
            15'b001001011001001 : data = 16'b1000111101010010;
            15'b001001011001010 : data = 16'b1000111100111110;
            15'b001001011001011 : data = 16'b1000111100101010;
            15'b001001011001100 : data = 16'b1000111100010101;
            15'b001001011001101 : data = 16'b1000111100000001;
            15'b001001011001110 : data = 16'b1000111011101100;
            15'b001001011001111 : data = 16'b1000111011011000;
            15'b001001011010000 : data = 16'b1000111011000011;
            15'b001001011010001 : data = 16'b1000111010101111;
            15'b001001011010010 : data = 16'b1000111010011010;
            15'b001001011010011 : data = 16'b1000111010000110;
            15'b001001011010100 : data = 16'b1000111001110001;
            15'b001001011010101 : data = 16'b1000111001011101;
            15'b001001011010110 : data = 16'b1000111001001001;
            15'b001001011010111 : data = 16'b1000111000110100;
            15'b001001011011000 : data = 16'b1000111000100000;
            15'b001001011011001 : data = 16'b1000111000001011;
            15'b001001011011010 : data = 16'b1000110111110111;
            15'b001001011011011 : data = 16'b1000110111100010;
            15'b001001011011100 : data = 16'b1000110111001110;
            15'b001001011011101 : data = 16'b1000110110111001;
            15'b001001011011110 : data = 16'b1000110110100101;
            15'b001001011011111 : data = 16'b1000110110010000;
            15'b001001011100000 : data = 16'b1000110101111100;
            15'b001001011100001 : data = 16'b1000110101100111;
            15'b001001011100010 : data = 16'b1000110101010011;
            15'b001001011100011 : data = 16'b1000110100111110;
            15'b001001011100100 : data = 16'b1000110100101010;
            15'b001001011100101 : data = 16'b1000110100010101;
            15'b001001011100110 : data = 16'b1000110100000001;
            15'b001001011100111 : data = 16'b1000110011101101;
            15'b001001011101000 : data = 16'b1000110011011000;
            15'b001001011101001 : data = 16'b1000110011000100;
            15'b001001011101010 : data = 16'b1000110010101111;
            15'b001001011101011 : data = 16'b1000110010011011;
            15'b001001011101100 : data = 16'b1000110010000110;
            15'b001001011101101 : data = 16'b1000110001110010;
            15'b001001011101110 : data = 16'b1000110001011101;
            15'b001001011101111 : data = 16'b1000110001001001;
            15'b001001011110000 : data = 16'b1000110000110100;
            15'b001001011110001 : data = 16'b1000110000100000;
            15'b001001011110010 : data = 16'b1000110000001011;
            15'b001001011110011 : data = 16'b1000101111110111;
            15'b001001011110100 : data = 16'b1000101111100010;
            15'b001001011110101 : data = 16'b1000101111001110;
            15'b001001011110110 : data = 16'b1000101110111001;
            15'b001001011110111 : data = 16'b1000101110100101;
            15'b001001011111000 : data = 16'b1000101110010000;
            15'b001001011111001 : data = 16'b1000101101111100;
            15'b001001011111010 : data = 16'b1000101101100111;
            15'b001001011111011 : data = 16'b1000101101010011;
            15'b001001011111100 : data = 16'b1000101100111110;
            15'b001001011111101 : data = 16'b1000101100101010;
            15'b001001011111110 : data = 16'b1000101100010101;
            15'b001001011111111 : data = 16'b1000101100000001;
            15'b001001100000000 : data = 16'b1000101011101100;
            15'b001001100000001 : data = 16'b1000101011011000;
            15'b001001100000010 : data = 16'b1000101011000011;
            15'b001001100000011 : data = 16'b1000101010101111;
            15'b001001100000100 : data = 16'b1000101010011010;
            15'b001001100000101 : data = 16'b1000101010000101;
            15'b001001100000110 : data = 16'b1000101001110001;
            15'b001001100000111 : data = 16'b1000101001011100;
            15'b001001100001000 : data = 16'b1000101001001000;
            15'b001001100001001 : data = 16'b1000101000110011;
            15'b001001100001010 : data = 16'b1000101000011111;
            15'b001001100001011 : data = 16'b1000101000001010;
            15'b001001100001100 : data = 16'b1000100111110110;
            15'b001001100001101 : data = 16'b1000100111100001;
            15'b001001100001110 : data = 16'b1000100111001101;
            15'b001001100001111 : data = 16'b1000100110111000;
            15'b001001100010000 : data = 16'b1000100110100100;
            15'b001001100010001 : data = 16'b1000100110001111;
            15'b001001100010010 : data = 16'b1000100101111011;
            15'b001001100010011 : data = 16'b1000100101100110;
            15'b001001100010100 : data = 16'b1000100101010010;
            15'b001001100010101 : data = 16'b1000100100111101;
            15'b001001100010110 : data = 16'b1000100100101001;
            15'b001001100010111 : data = 16'b1000100100010100;
            15'b001001100011000 : data = 16'b1000100011111111;
            15'b001001100011001 : data = 16'b1000100011101011;
            15'b001001100011010 : data = 16'b1000100011010110;
            15'b001001100011011 : data = 16'b1000100011000010;
            15'b001001100011100 : data = 16'b1000100010101101;
            15'b001001100011101 : data = 16'b1000100010011001;
            15'b001001100011110 : data = 16'b1000100010000100;
            15'b001001100011111 : data = 16'b1000100001110000;
            15'b001001100100000 : data = 16'b1000100001011011;
            15'b001001100100001 : data = 16'b1000100001000111;
            15'b001001100100010 : data = 16'b1000100000110010;
            15'b001001100100011 : data = 16'b1000100000011110;
            15'b001001100100100 : data = 16'b1000100000001001;
            15'b001001100100101 : data = 16'b1000011111110100;
            15'b001001100100110 : data = 16'b1000011111100000;
            15'b001001100100111 : data = 16'b1000011111001011;
            15'b001001100101000 : data = 16'b1000011110110111;
            15'b001001100101001 : data = 16'b1000011110100010;
            15'b001001100101010 : data = 16'b1000011110001110;
            15'b001001100101011 : data = 16'b1000011101111001;
            15'b001001100101100 : data = 16'b1000011101100101;
            15'b001001100101101 : data = 16'b1000011101010000;
            15'b001001100101110 : data = 16'b1000011100111011;
            15'b001001100101111 : data = 16'b1000011100100111;
            15'b001001100110000 : data = 16'b1000011100010010;
            15'b001001100110001 : data = 16'b1000011011111110;
            15'b001001100110010 : data = 16'b1000011011101001;
            15'b001001100110011 : data = 16'b1000011011010101;
            15'b001001100110100 : data = 16'b1000011011000000;
            15'b001001100110101 : data = 16'b1000011010101100;
            15'b001001100110110 : data = 16'b1000011010010111;
            15'b001001100110111 : data = 16'b1000011010000010;
            15'b001001100111000 : data = 16'b1000011001101110;
            15'b001001100111001 : data = 16'b1000011001011001;
            15'b001001100111010 : data = 16'b1000011001000101;
            15'b001001100111011 : data = 16'b1000011000110000;
            15'b001001100111100 : data = 16'b1000011000011100;
            15'b001001100111101 : data = 16'b1000011000000111;
            15'b001001100111110 : data = 16'b1000010111110010;
            15'b001001100111111 : data = 16'b1000010111011110;
            15'b001001101000000 : data = 16'b1000010111001001;
            15'b001001101000001 : data = 16'b1000010110110101;
            15'b001001101000010 : data = 16'b1000010110100000;
            15'b001001101000011 : data = 16'b1000010110001100;
            15'b001001101000100 : data = 16'b1000010101110111;
            15'b001001101000101 : data = 16'b1000010101100010;
            15'b001001101000110 : data = 16'b1000010101001110;
            15'b001001101000111 : data = 16'b1000010100111001;
            15'b001001101001000 : data = 16'b1000010100100101;
            15'b001001101001001 : data = 16'b1000010100010000;
            15'b001001101001010 : data = 16'b1000010011111100;
            15'b001001101001011 : data = 16'b1000010011100111;
            15'b001001101001100 : data = 16'b1000010011010010;
            15'b001001101001101 : data = 16'b1000010010111110;
            15'b001001101001110 : data = 16'b1000010010101001;
            15'b001001101001111 : data = 16'b1000010010010101;
            15'b001001101010000 : data = 16'b1000010010000000;
            15'b001001101010001 : data = 16'b1000010001101100;
            15'b001001101010010 : data = 16'b1000010001010111;
            15'b001001101010011 : data = 16'b1000010001000010;
            15'b001001101010100 : data = 16'b1000010000101110;
            15'b001001101010101 : data = 16'b1000010000011001;
            15'b001001101010110 : data = 16'b1000010000000101;
            15'b001001101010111 : data = 16'b1000001111110000;
            15'b001001101011000 : data = 16'b1000001111011100;
            15'b001001101011001 : data = 16'b1000001111000111;
            15'b001001101011010 : data = 16'b1000001110110010;
            15'b001001101011011 : data = 16'b1000001110011110;
            15'b001001101011100 : data = 16'b1000001110001001;
            15'b001001101011101 : data = 16'b1000001101110101;
            15'b001001101011110 : data = 16'b1000001101100000;
            15'b001001101011111 : data = 16'b1000001101001100;
            15'b001001101100000 : data = 16'b1000001100110111;
            15'b001001101100001 : data = 16'b1000001100100010;
            15'b001001101100010 : data = 16'b1000001100001110;
            15'b001001101100011 : data = 16'b1000001011111001;
            15'b001001101100100 : data = 16'b1000001011100101;
            15'b001001101100101 : data = 16'b1000001011010000;
            15'b001001101100110 : data = 16'b1000001010111011;
            15'b001001101100111 : data = 16'b1000001010100111;
            15'b001001101101000 : data = 16'b1000001010010010;
            15'b001001101101001 : data = 16'b1000001001111110;
            15'b001001101101010 : data = 16'b1000001001101001;
            15'b001001101101011 : data = 16'b1000001001010101;
            15'b001001101101100 : data = 16'b1000001001000000;
            15'b001001101101101 : data = 16'b1000001000101011;
            15'b001001101101110 : data = 16'b1000001000010111;
            15'b001001101101111 : data = 16'b1000001000000010;
            15'b001001101110000 : data = 16'b1000000111101110;
            15'b001001101110001 : data = 16'b1000000111011001;
            15'b001001101110010 : data = 16'b1000000111000100;
            15'b001001101110011 : data = 16'b1000000110110000;
            15'b001001101110100 : data = 16'b1000000110011011;
            15'b001001101110101 : data = 16'b1000000110000111;
            15'b001001101110110 : data = 16'b1000000101110010;
            15'b001001101110111 : data = 16'b1000000101011101;
            15'b001001101111000 : data = 16'b1000000101001001;
            15'b001001101111001 : data = 16'b1000000100110100;
            15'b001001101111010 : data = 16'b1000000100100000;
            15'b001001101111011 : data = 16'b1000000100001011;
            15'b001001101111100 : data = 16'b1000000011110111;
            15'b001001101111101 : data = 16'b1000000011100010;
            15'b001001101111110 : data = 16'b1000000011001101;
            15'b001001101111111 : data = 16'b1000000010111001;
            15'b001001110000000 : data = 16'b1000000010100100;
            15'b001001110000001 : data = 16'b1000000010010000;
            15'b001001110000010 : data = 16'b1000000001111011;
            15'b001001110000011 : data = 16'b1000000001100110;
            15'b001001110000100 : data = 16'b1000000001010010;
            15'b001001110000101 : data = 16'b1000000000111101;
            15'b001001110000110 : data = 16'b1000000000101001;
            15'b001001110000111 : data = 16'b1000000000010100;
            15'b001001110001000 : data = 16'b1000000000000000;
            15'b001001110001001 : data = 16'b0111111111101011;
            15'b001001110001010 : data = 16'b0111111111010110;
            15'b001001110001011 : data = 16'b0111111111000010;
            15'b001001110001100 : data = 16'b0111111110101101;
            15'b001001110001101 : data = 16'b0111111110011001;
            15'b001001110001110 : data = 16'b0111111110000100;
            15'b001001110001111 : data = 16'b0111111101101111;
            15'b001001110010000 : data = 16'b0111111101011011;
            15'b001001110010001 : data = 16'b0111111101000110;
            15'b001001110010010 : data = 16'b0111111100110010;
            15'b001001110010011 : data = 16'b0111111100011101;
            15'b001001110010100 : data = 16'b0111111100001000;
            15'b001001110010101 : data = 16'b0111111011110100;
            15'b001001110010110 : data = 16'b0111111011011111;
            15'b001001110010111 : data = 16'b0111111011001011;
            15'b001001110011000 : data = 16'b0111111010110110;
            15'b001001110011001 : data = 16'b0111111010100010;
            15'b001001110011010 : data = 16'b0111111010001101;
            15'b001001110011011 : data = 16'b0111111001111000;
            15'b001001110011100 : data = 16'b0111111001100100;
            15'b001001110011101 : data = 16'b0111111001001111;
            15'b001001110011110 : data = 16'b0111111000111011;
            15'b001001110011111 : data = 16'b0111111000100110;
            15'b001001110100000 : data = 16'b0111111000010001;
            15'b001001110100001 : data = 16'b0111110111111101;
            15'b001001110100010 : data = 16'b0111110111101000;
            15'b001001110100011 : data = 16'b0111110111010100;
            15'b001001110100100 : data = 16'b0111110110111111;
            15'b001001110100101 : data = 16'b0111110110101010;
            15'b001001110100110 : data = 16'b0111110110010110;
            15'b001001110100111 : data = 16'b0111110110000001;
            15'b001001110101000 : data = 16'b0111110101101101;
            15'b001001110101001 : data = 16'b0111110101011000;
            15'b001001110101010 : data = 16'b0111110101000100;
            15'b001001110101011 : data = 16'b0111110100101111;
            15'b001001110101100 : data = 16'b0111110100011010;
            15'b001001110101101 : data = 16'b0111110100000110;
            15'b001001110101110 : data = 16'b0111110011110001;
            15'b001001110101111 : data = 16'b0111110011011101;
            15'b001001110110000 : data = 16'b0111110011001000;
            15'b001001110110001 : data = 16'b0111110010110011;
            15'b001001110110010 : data = 16'b0111110010011111;
            15'b001001110110011 : data = 16'b0111110010001010;
            15'b001001110110100 : data = 16'b0111110001110110;
            15'b001001110110101 : data = 16'b0111110001100001;
            15'b001001110110110 : data = 16'b0111110001001101;
            15'b001001110110111 : data = 16'b0111110000111000;
            15'b001001110111000 : data = 16'b0111110000100011;
            15'b001001110111001 : data = 16'b0111110000001111;
            15'b001001110111010 : data = 16'b0111101111111010;
            15'b001001110111011 : data = 16'b0111101111100110;
            15'b001001110111100 : data = 16'b0111101111010001;
            15'b001001110111101 : data = 16'b0111101110111101;
            15'b001001110111110 : data = 16'b0111101110101000;
            15'b001001110111111 : data = 16'b0111101110010011;
            15'b001001111000000 : data = 16'b0111101101111111;
            15'b001001111000001 : data = 16'b0111101101101010;
            15'b001001111000010 : data = 16'b0111101101010110;
            15'b001001111000011 : data = 16'b0111101101000001;
            15'b001001111000100 : data = 16'b0111101100101101;
            15'b001001111000101 : data = 16'b0111101100011000;
            15'b001001111000110 : data = 16'b0111101100000011;
            15'b001001111000111 : data = 16'b0111101011101111;
            15'b001001111001000 : data = 16'b0111101011011010;
            15'b001001111001001 : data = 16'b0111101011000110;
            15'b001001111001010 : data = 16'b0111101010110001;
            15'b001001111001011 : data = 16'b0111101010011101;
            15'b001001111001100 : data = 16'b0111101010001000;
            15'b001001111001101 : data = 16'b0111101001110011;
            15'b001001111001110 : data = 16'b0111101001011111;
            15'b001001111001111 : data = 16'b0111101001001010;
            15'b001001111010000 : data = 16'b0111101000110110;
            15'b001001111010001 : data = 16'b0111101000100001;
            15'b001001111010010 : data = 16'b0111101000001101;
            15'b001001111010011 : data = 16'b0111100111111000;
            15'b001001111010100 : data = 16'b0111100111100011;
            15'b001001111010101 : data = 16'b0111100111001111;
            15'b001001111010110 : data = 16'b0111100110111010;
            15'b001001111010111 : data = 16'b0111100110100110;
            15'b001001111011000 : data = 16'b0111100110010001;
            15'b001001111011001 : data = 16'b0111100101111101;
            15'b001001111011010 : data = 16'b0111100101101000;
            15'b001001111011011 : data = 16'b0111100101010011;
            15'b001001111011100 : data = 16'b0111100100111111;
            15'b001001111011101 : data = 16'b0111100100101010;
            15'b001001111011110 : data = 16'b0111100100010110;
            15'b001001111011111 : data = 16'b0111100100000001;
            15'b001001111100000 : data = 16'b0111100011101101;
            15'b001001111100001 : data = 16'b0111100011011000;
            15'b001001111100010 : data = 16'b0111100011000100;
            15'b001001111100011 : data = 16'b0111100010101111;
            15'b001001111100100 : data = 16'b0111100010011010;
            15'b001001111100101 : data = 16'b0111100010000110;
            15'b001001111100110 : data = 16'b0111100001110001;
            15'b001001111100111 : data = 16'b0111100001011101;
            15'b001001111101000 : data = 16'b0111100001001000;
            15'b001001111101001 : data = 16'b0111100000110100;
            15'b001001111101010 : data = 16'b0111100000011111;
            15'b001001111101011 : data = 16'b0111100000001011;
            15'b001001111101100 : data = 16'b0111011111110110;
            15'b001001111101101 : data = 16'b0111011111100001;
            15'b001001111101110 : data = 16'b0111011111001101;
            15'b001001111101111 : data = 16'b0111011110111000;
            15'b001001111110000 : data = 16'b0111011110100100;
            15'b001001111110001 : data = 16'b0111011110001111;
            15'b001001111110010 : data = 16'b0111011101111011;
            15'b001001111110011 : data = 16'b0111011101100110;
            15'b001001111110100 : data = 16'b0111011101010010;
            15'b001001111110101 : data = 16'b0111011100111101;
            15'b001001111110110 : data = 16'b0111011100101001;
            15'b001001111110111 : data = 16'b0111011100010100;
            15'b001001111111000 : data = 16'b0111011100000000;
            15'b001001111111001 : data = 16'b0111011011101011;
            15'b001001111111010 : data = 16'b0111011011010110;
            15'b001001111111011 : data = 16'b0111011011000010;
            15'b001001111111100 : data = 16'b0111011010101101;
            15'b001001111111101 : data = 16'b0111011010011001;
            15'b001001111111110 : data = 16'b0111011010000100;
            15'b001001111111111 : data = 16'b0111011001110000;
            15'b001010000000000 : data = 16'b0111011001011011;
            15'b001010000000001 : data = 16'b0111011001000111;
            15'b001010000000010 : data = 16'b0111011000110010;
            15'b001010000000011 : data = 16'b0111011000011110;
            15'b001010000000100 : data = 16'b0111011000001001;
            15'b001010000000101 : data = 16'b0111010111110101;
            15'b001010000000110 : data = 16'b0111010111100000;
            15'b001010000000111 : data = 16'b0111010111001100;
            15'b001010000001000 : data = 16'b0111010110110111;
            15'b001010000001001 : data = 16'b0111010110100011;
            15'b001010000001010 : data = 16'b0111010110001110;
            15'b001010000001011 : data = 16'b0111010101111010;
            15'b001010000001100 : data = 16'b0111010101100101;
            15'b001010000001101 : data = 16'b0111010101010000;
            15'b001010000001110 : data = 16'b0111010100111100;
            15'b001010000001111 : data = 16'b0111010100100111;
            15'b001010000010000 : data = 16'b0111010100010011;
            15'b001010000010001 : data = 16'b0111010011111110;
            15'b001010000010010 : data = 16'b0111010011101010;
            15'b001010000010011 : data = 16'b0111010011010101;
            15'b001010000010100 : data = 16'b0111010011000001;
            15'b001010000010101 : data = 16'b0111010010101100;
            15'b001010000010110 : data = 16'b0111010010011000;
            15'b001010000010111 : data = 16'b0111010010000011;
            15'b001010000011000 : data = 16'b0111010001101111;
            15'b001010000011001 : data = 16'b0111010001011010;
            15'b001010000011010 : data = 16'b0111010001000110;
            15'b001010000011011 : data = 16'b0111010000110001;
            15'b001010000011100 : data = 16'b0111010000011101;
            15'b001010000011101 : data = 16'b0111010000001000;
            15'b001010000011110 : data = 16'b0111001111110100;
            15'b001010000011111 : data = 16'b0111001111011111;
            15'b001010000100000 : data = 16'b0111001111001011;
            15'b001010000100001 : data = 16'b0111001110110110;
            15'b001010000100010 : data = 16'b0111001110100010;
            15'b001010000100011 : data = 16'b0111001110001101;
            15'b001010000100100 : data = 16'b0111001101111001;
            15'b001010000100101 : data = 16'b0111001101100100;
            15'b001010000100110 : data = 16'b0111001101010000;
            15'b001010000100111 : data = 16'b0111001100111011;
            15'b001010000101000 : data = 16'b0111001100100111;
            15'b001010000101001 : data = 16'b0111001100010010;
            15'b001010000101010 : data = 16'b0111001011111110;
            15'b001010000101011 : data = 16'b0111001011101010;
            15'b001010000101100 : data = 16'b0111001011010101;
            15'b001010000101101 : data = 16'b0111001011000001;
            15'b001010000101110 : data = 16'b0111001010101100;
            15'b001010000101111 : data = 16'b0111001010011000;
            15'b001010000110000 : data = 16'b0111001010000011;
            15'b001010000110001 : data = 16'b0111001001101111;
            15'b001010000110010 : data = 16'b0111001001011010;
            15'b001010000110011 : data = 16'b0111001001000110;
            15'b001010000110100 : data = 16'b0111001000110001;
            15'b001010000110101 : data = 16'b0111001000011101;
            15'b001010000110110 : data = 16'b0111001000001000;
            15'b001010000110111 : data = 16'b0111000111110100;
            15'b001010000111000 : data = 16'b0111000111011111;
            15'b001010000111001 : data = 16'b0111000111001011;
            15'b001010000111010 : data = 16'b0111000110110110;
            15'b001010000111011 : data = 16'b0111000110100010;
            15'b001010000111100 : data = 16'b0111000110001110;
            15'b001010000111101 : data = 16'b0111000101111001;
            15'b001010000111110 : data = 16'b0111000101100101;
            15'b001010000111111 : data = 16'b0111000101010000;
            15'b001010001000000 : data = 16'b0111000100111100;
            15'b001010001000001 : data = 16'b0111000100100111;
            15'b001010001000010 : data = 16'b0111000100010011;
            15'b001010001000011 : data = 16'b0111000011111110;
            15'b001010001000100 : data = 16'b0111000011101010;
            15'b001010001000101 : data = 16'b0111000011010101;
            15'b001010001000110 : data = 16'b0111000011000001;
            15'b001010001000111 : data = 16'b0111000010101101;
            15'b001010001001000 : data = 16'b0111000010011000;
            15'b001010001001001 : data = 16'b0111000010000100;
            15'b001010001001010 : data = 16'b0111000001101111;
            15'b001010001001011 : data = 16'b0111000001011011;
            15'b001010001001100 : data = 16'b0111000001000110;
            15'b001010001001101 : data = 16'b0111000000110010;
            15'b001010001001110 : data = 16'b0111000000011110;
            15'b001010001001111 : data = 16'b0111000000001001;
            15'b001010001010000 : data = 16'b0110111111110101;
            15'b001010001010001 : data = 16'b0110111111100000;
            15'b001010001010010 : data = 16'b0110111111001100;
            15'b001010001010011 : data = 16'b0110111110110111;
            15'b001010001010100 : data = 16'b0110111110100011;
            15'b001010001010101 : data = 16'b0110111110001111;
            15'b001010001010110 : data = 16'b0110111101111010;
            15'b001010001010111 : data = 16'b0110111101100110;
            15'b001010001011000 : data = 16'b0110111101010001;
            15'b001010001011001 : data = 16'b0110111100111101;
            15'b001010001011010 : data = 16'b0110111100101001;
            15'b001010001011011 : data = 16'b0110111100010100;
            15'b001010001011100 : data = 16'b0110111100000000;
            15'b001010001011101 : data = 16'b0110111011101011;
            15'b001010001011110 : data = 16'b0110111011010111;
            15'b001010001011111 : data = 16'b0110111011000011;
            15'b001010001100000 : data = 16'b0110111010101110;
            15'b001010001100001 : data = 16'b0110111010011010;
            15'b001010001100010 : data = 16'b0110111010000101;
            15'b001010001100011 : data = 16'b0110111001110001;
            15'b001010001100100 : data = 16'b0110111001011101;
            15'b001010001100101 : data = 16'b0110111001001000;
            15'b001010001100110 : data = 16'b0110111000110100;
            15'b001010001100111 : data = 16'b0110111000011111;
            15'b001010001101000 : data = 16'b0110111000001011;
            15'b001010001101001 : data = 16'b0110110111110111;
            15'b001010001101010 : data = 16'b0110110111100010;
            15'b001010001101011 : data = 16'b0110110111001110;
            15'b001010001101100 : data = 16'b0110110110111001;
            15'b001010001101101 : data = 16'b0110110110100101;
            15'b001010001101110 : data = 16'b0110110110010001;
            15'b001010001101111 : data = 16'b0110110101111100;
            15'b001010001110000 : data = 16'b0110110101101000;
            15'b001010001110001 : data = 16'b0110110101010100;
            15'b001010001110010 : data = 16'b0110110100111111;
            15'b001010001110011 : data = 16'b0110110100101011;
            15'b001010001110100 : data = 16'b0110110100010110;
            15'b001010001110101 : data = 16'b0110110100000010;
            15'b001010001110110 : data = 16'b0110110011101110;
            15'b001010001110111 : data = 16'b0110110011011001;
            15'b001010001111000 : data = 16'b0110110011000101;
            15'b001010001111001 : data = 16'b0110110010110001;
            15'b001010001111010 : data = 16'b0110110010011100;
            15'b001010001111011 : data = 16'b0110110010001000;
            15'b001010001111100 : data = 16'b0110110001110100;
            15'b001010001111101 : data = 16'b0110110001011111;
            15'b001010001111110 : data = 16'b0110110001001011;
            15'b001010001111111 : data = 16'b0110110000110111;
            15'b001010010000000 : data = 16'b0110110000100010;
            15'b001010010000001 : data = 16'b0110110000001110;
            15'b001010010000010 : data = 16'b0110101111111010;
            15'b001010010000011 : data = 16'b0110101111100101;
            15'b001010010000100 : data = 16'b0110101111010001;
            15'b001010010000101 : data = 16'b0110101110111101;
            15'b001010010000110 : data = 16'b0110101110101000;
            15'b001010010000111 : data = 16'b0110101110010100;
            15'b001010010001000 : data = 16'b0110101110000000;
            15'b001010010001001 : data = 16'b0110101101101011;
            15'b001010010001010 : data = 16'b0110101101010111;
            15'b001010010001011 : data = 16'b0110101101000011;
            15'b001010010001100 : data = 16'b0110101100101110;
            15'b001010010001101 : data = 16'b0110101100011010;
            15'b001010010001110 : data = 16'b0110101100000110;
            15'b001010010001111 : data = 16'b0110101011110001;
            15'b001010010010000 : data = 16'b0110101011011101;
            15'b001010010010001 : data = 16'b0110101011001001;
            15'b001010010010010 : data = 16'b0110101010110101;
            15'b001010010010011 : data = 16'b0110101010100000;
            15'b001010010010100 : data = 16'b0110101010001100;
            15'b001010010010101 : data = 16'b0110101001111000;
            15'b001010010010110 : data = 16'b0110101001100011;
            15'b001010010010111 : data = 16'b0110101001001111;
            15'b001010010011000 : data = 16'b0110101000111011;
            15'b001010010011001 : data = 16'b0110101000100110;
            15'b001010010011010 : data = 16'b0110101000010010;
            15'b001010010011011 : data = 16'b0110100111111110;
            15'b001010010011100 : data = 16'b0110100111101010;
            15'b001010010011101 : data = 16'b0110100111010101;
            15'b001010010011110 : data = 16'b0110100111000001;
            15'b001010010011111 : data = 16'b0110100110101101;
            15'b001010010100000 : data = 16'b0110100110011001;
            15'b001010010100001 : data = 16'b0110100110000100;
            15'b001010010100010 : data = 16'b0110100101110000;
            15'b001010010100011 : data = 16'b0110100101011100;
            15'b001010010100100 : data = 16'b0110100101000111;
            15'b001010010100101 : data = 16'b0110100100110011;
            15'b001010010100110 : data = 16'b0110100100011111;
            15'b001010010100111 : data = 16'b0110100100001011;
            15'b001010010101000 : data = 16'b0110100011110110;
            15'b001010010101001 : data = 16'b0110100011100010;
            15'b001010010101010 : data = 16'b0110100011001110;
            15'b001010010101011 : data = 16'b0110100010111010;
            15'b001010010101100 : data = 16'b0110100010100101;
            15'b001010010101101 : data = 16'b0110100010010001;
            15'b001010010101110 : data = 16'b0110100001111101;
            15'b001010010101111 : data = 16'b0110100001101001;
            15'b001010010110000 : data = 16'b0110100001010100;
            15'b001010010110001 : data = 16'b0110100001000000;
            15'b001010010110010 : data = 16'b0110100000101100;
            15'b001010010110011 : data = 16'b0110100000011000;
            15'b001010010110100 : data = 16'b0110100000000100;
            15'b001010010110101 : data = 16'b0110011111101111;
            15'b001010010110110 : data = 16'b0110011111011011;
            15'b001010010110111 : data = 16'b0110011111000111;
            15'b001010010111000 : data = 16'b0110011110110011;
            15'b001010010111001 : data = 16'b0110011110011110;
            15'b001010010111010 : data = 16'b0110011110001010;
            15'b001010010111011 : data = 16'b0110011101110110;
            15'b001010010111100 : data = 16'b0110011101100010;
            15'b001010010111101 : data = 16'b0110011101001110;
            15'b001010010111110 : data = 16'b0110011100111001;
            15'b001010010111111 : data = 16'b0110011100100101;
            15'b001010011000000 : data = 16'b0110011100010001;
            15'b001010011000001 : data = 16'b0110011011111101;
            15'b001010011000010 : data = 16'b0110011011101001;
            15'b001010011000011 : data = 16'b0110011011010101;
            15'b001010011000100 : data = 16'b0110011011000000;
            15'b001010011000101 : data = 16'b0110011010101100;
            15'b001010011000110 : data = 16'b0110011010011000;
            15'b001010011000111 : data = 16'b0110011010000100;
            15'b001010011001000 : data = 16'b0110011001110000;
            15'b001010011001001 : data = 16'b0110011001011011;
            15'b001010011001010 : data = 16'b0110011001000111;
            15'b001010011001011 : data = 16'b0110011000110011;
            15'b001010011001100 : data = 16'b0110011000011111;
            15'b001010011001101 : data = 16'b0110011000001011;
            15'b001010011001110 : data = 16'b0110010111110111;
            15'b001010011001111 : data = 16'b0110010111100010;
            15'b001010011010000 : data = 16'b0110010111001110;
            15'b001010011010001 : data = 16'b0110010110111010;
            15'b001010011010010 : data = 16'b0110010110100110;
            15'b001010011010011 : data = 16'b0110010110010010;
            15'b001010011010100 : data = 16'b0110010101111110;
            15'b001010011010101 : data = 16'b0110010101101010;
            15'b001010011010110 : data = 16'b0110010101010101;
            15'b001010011010111 : data = 16'b0110010101000001;
            15'b001010011011000 : data = 16'b0110010100101101;
            15'b001010011011001 : data = 16'b0110010100011001;
            15'b001010011011010 : data = 16'b0110010100000101;
            15'b001010011011011 : data = 16'b0110010011110001;
            15'b001010011011100 : data = 16'b0110010011011101;
            15'b001010011011101 : data = 16'b0110010011001001;
            15'b001010011011110 : data = 16'b0110010010110100;
            15'b001010011011111 : data = 16'b0110010010100000;
            15'b001010011100000 : data = 16'b0110010010001100;
            15'b001010011100001 : data = 16'b0110010001111000;
            15'b001010011100010 : data = 16'b0110010001100100;
            15'b001010011100011 : data = 16'b0110010001010000;
            15'b001010011100100 : data = 16'b0110010000111100;
            15'b001010011100101 : data = 16'b0110010000101000;
            15'b001010011100110 : data = 16'b0110010000010100;
            15'b001010011100111 : data = 16'b0110010000000000;
            15'b001010011101000 : data = 16'b0110001111101011;
            15'b001010011101001 : data = 16'b0110001111010111;
            15'b001010011101010 : data = 16'b0110001111000011;
            15'b001010011101011 : data = 16'b0110001110101111;
            15'b001010011101100 : data = 16'b0110001110011011;
            15'b001010011101101 : data = 16'b0110001110000111;
            15'b001010011101110 : data = 16'b0110001101110011;
            15'b001010011101111 : data = 16'b0110001101011111;
            15'b001010011110000 : data = 16'b0110001101001011;
            15'b001010011110001 : data = 16'b0110001100110111;
            15'b001010011110010 : data = 16'b0110001100100011;
            15'b001010011110011 : data = 16'b0110001100001111;
            15'b001010011110100 : data = 16'b0110001011111011;
            15'b001010011110101 : data = 16'b0110001011100111;
            15'b001010011110110 : data = 16'b0110001011010010;
            15'b001010011110111 : data = 16'b0110001010111110;
            15'b001010011111000 : data = 16'b0110001010101010;
            15'b001010011111001 : data = 16'b0110001010010110;
            15'b001010011111010 : data = 16'b0110001010000010;
            15'b001010011111011 : data = 16'b0110001001101110;
            15'b001010011111100 : data = 16'b0110001001011010;
            15'b001010011111101 : data = 16'b0110001001000110;
            15'b001010011111110 : data = 16'b0110001000110010;
            15'b001010011111111 : data = 16'b0110001000011110;
            15'b001010100000000 : data = 16'b0110001000001010;
            15'b001010100000001 : data = 16'b0110000111110110;
            15'b001010100000010 : data = 16'b0110000111100010;
            15'b001010100000011 : data = 16'b0110000111001110;
            15'b001010100000100 : data = 16'b0110000110111010;
            15'b001010100000101 : data = 16'b0110000110100110;
            15'b001010100000110 : data = 16'b0110000110010010;
            15'b001010100000111 : data = 16'b0110000101111110;
            15'b001010100001000 : data = 16'b0110000101101010;
            15'b001010100001001 : data = 16'b0110000101010110;
            15'b001010100001010 : data = 16'b0110000101000010;
            15'b001010100001011 : data = 16'b0110000100101110;
            15'b001010100001100 : data = 16'b0110000100011010;
            15'b001010100001101 : data = 16'b0110000100000110;
            15'b001010100001110 : data = 16'b0110000011110010;
            15'b001010100001111 : data = 16'b0110000011011110;
            15'b001010100010000 : data = 16'b0110000011001010;
            15'b001010100010001 : data = 16'b0110000010110110;
            15'b001010100010010 : data = 16'b0110000010100010;
            15'b001010100010011 : data = 16'b0110000010001110;
            15'b001010100010100 : data = 16'b0110000001111010;
            15'b001010100010101 : data = 16'b0110000001100111;
            15'b001010100010110 : data = 16'b0110000001010011;
            15'b001010100010111 : data = 16'b0110000000111111;
            15'b001010100011000 : data = 16'b0110000000101011;
            15'b001010100011001 : data = 16'b0110000000010111;
            15'b001010100011010 : data = 16'b0110000000000011;
            15'b001010100011011 : data = 16'b0101111111101111;
            15'b001010100011100 : data = 16'b0101111111011011;
            15'b001010100011101 : data = 16'b0101111111000111;
            15'b001010100011110 : data = 16'b0101111110110011;
            15'b001010100011111 : data = 16'b0101111110011111;
            15'b001010100100000 : data = 16'b0101111110001011;
            15'b001010100100001 : data = 16'b0101111101110111;
            15'b001010100100010 : data = 16'b0101111101100011;
            15'b001010100100011 : data = 16'b0101111101010000;
            15'b001010100100100 : data = 16'b0101111100111100;
            15'b001010100100101 : data = 16'b0101111100101000;
            15'b001010100100110 : data = 16'b0101111100010100;
            15'b001010100100111 : data = 16'b0101111100000000;
            15'b001010100101000 : data = 16'b0101111011101100;
            15'b001010100101001 : data = 16'b0101111011011000;
            15'b001010100101010 : data = 16'b0101111011000100;
            15'b001010100101011 : data = 16'b0101111010110000;
            15'b001010100101100 : data = 16'b0101111010011101;
            15'b001010100101101 : data = 16'b0101111010001001;
            15'b001010100101110 : data = 16'b0101111001110101;
            15'b001010100101111 : data = 16'b0101111001100001;
            15'b001010100110000 : data = 16'b0101111001001101;
            15'b001010100110001 : data = 16'b0101111000111001;
            15'b001010100110010 : data = 16'b0101111000100101;
            15'b001010100110011 : data = 16'b0101111000010001;
            15'b001010100110100 : data = 16'b0101110111111110;
            15'b001010100110101 : data = 16'b0101110111101010;
            15'b001010100110110 : data = 16'b0101110111010110;
            15'b001010100110111 : data = 16'b0101110111000010;
            15'b001010100111000 : data = 16'b0101110110101110;
            15'b001010100111001 : data = 16'b0101110110011010;
            15'b001010100111010 : data = 16'b0101110110000111;
            15'b001010100111011 : data = 16'b0101110101110011;
            15'b001010100111100 : data = 16'b0101110101011111;
            15'b001010100111101 : data = 16'b0101110101001011;
            15'b001010100111110 : data = 16'b0101110100110111;
            15'b001010100111111 : data = 16'b0101110100100011;
            15'b001010101000000 : data = 16'b0101110100010000;
            15'b001010101000001 : data = 16'b0101110011111100;
            15'b001010101000010 : data = 16'b0101110011101000;
            15'b001010101000011 : data = 16'b0101110011010100;
            15'b001010101000100 : data = 16'b0101110011000000;
            15'b001010101000101 : data = 16'b0101110010101101;
            15'b001010101000110 : data = 16'b0101110010011001;
            15'b001010101000111 : data = 16'b0101110010000101;
            15'b001010101001000 : data = 16'b0101110001110001;
            15'b001010101001001 : data = 16'b0101110001011110;
            15'b001010101001010 : data = 16'b0101110001001010;
            15'b001010101001011 : data = 16'b0101110000110110;
            15'b001010101001100 : data = 16'b0101110000100010;
            15'b001010101001101 : data = 16'b0101110000001111;
            15'b001010101001110 : data = 16'b0101101111111011;
            15'b001010101001111 : data = 16'b0101101111100111;
            15'b001010101010000 : data = 16'b0101101111010011;
            15'b001010101010001 : data = 16'b0101101110111111;
            15'b001010101010010 : data = 16'b0101101110101100;
            15'b001010101010011 : data = 16'b0101101110011000;
            15'b001010101010100 : data = 16'b0101101110000100;
            15'b001010101010101 : data = 16'b0101101101110001;
            15'b001010101010110 : data = 16'b0101101101011101;
            15'b001010101010111 : data = 16'b0101101101001001;
            15'b001010101011000 : data = 16'b0101101100110101;
            15'b001010101011001 : data = 16'b0101101100100010;
            15'b001010101011010 : data = 16'b0101101100001110;
            15'b001010101011011 : data = 16'b0101101011111010;
            15'b001010101011100 : data = 16'b0101101011100111;
            15'b001010101011101 : data = 16'b0101101011010011;
            15'b001010101011110 : data = 16'b0101101010111111;
            15'b001010101011111 : data = 16'b0101101010101011;
            15'b001010101100000 : data = 16'b0101101010011000;
            15'b001010101100001 : data = 16'b0101101010000100;
            15'b001010101100010 : data = 16'b0101101001110000;
            15'b001010101100011 : data = 16'b0101101001011101;
            15'b001010101100100 : data = 16'b0101101001001001;
            15'b001010101100101 : data = 16'b0101101000110101;
            15'b001010101100110 : data = 16'b0101101000100010;
            15'b001010101100111 : data = 16'b0101101000001110;
            15'b001010101101000 : data = 16'b0101100111111010;
            15'b001010101101001 : data = 16'b0101100111100111;
            15'b001010101101010 : data = 16'b0101100111010011;
            15'b001010101101011 : data = 16'b0101100110111111;
            15'b001010101101100 : data = 16'b0101100110101100;
            15'b001010101101101 : data = 16'b0101100110011000;
            15'b001010101101110 : data = 16'b0101100110000100;
            15'b001010101101111 : data = 16'b0101100101110001;
            15'b001010101110000 : data = 16'b0101100101011101;
            15'b001010101110001 : data = 16'b0101100101001010;
            15'b001010101110010 : data = 16'b0101100100110110;
            15'b001010101110011 : data = 16'b0101100100100010;
            15'b001010101110100 : data = 16'b0101100100001111;
            15'b001010101110101 : data = 16'b0101100011111011;
            15'b001010101110110 : data = 16'b0101100011100111;
            15'b001010101110111 : data = 16'b0101100011010100;
            15'b001010101111000 : data = 16'b0101100011000000;
            15'b001010101111001 : data = 16'b0101100010101101;
            15'b001010101111010 : data = 16'b0101100010011001;
            15'b001010101111011 : data = 16'b0101100010000110;
            15'b001010101111100 : data = 16'b0101100001110010;
            15'b001010101111101 : data = 16'b0101100001011110;
            15'b001010101111110 : data = 16'b0101100001001011;
            15'b001010101111111 : data = 16'b0101100000110111;
            15'b001010110000000 : data = 16'b0101100000100100;
            15'b001010110000001 : data = 16'b0101100000010000;
            15'b001010110000010 : data = 16'b0101011111111101;
            15'b001010110000011 : data = 16'b0101011111101001;
            15'b001010110000100 : data = 16'b0101011111010101;
            15'b001010110000101 : data = 16'b0101011111000010;
            15'b001010110000110 : data = 16'b0101011110101110;
            15'b001010110000111 : data = 16'b0101011110011011;
            15'b001010110001000 : data = 16'b0101011110000111;
            15'b001010110001001 : data = 16'b0101011101110100;
            15'b001010110001010 : data = 16'b0101011101100000;
            15'b001010110001011 : data = 16'b0101011101001101;
            15'b001010110001100 : data = 16'b0101011100111001;
            15'b001010110001101 : data = 16'b0101011100100110;
            15'b001010110001110 : data = 16'b0101011100010010;
            15'b001010110001111 : data = 16'b0101011011111111;
            15'b001010110010000 : data = 16'b0101011011101011;
            15'b001010110010001 : data = 16'b0101011011011000;
            15'b001010110010010 : data = 16'b0101011011000100;
            15'b001010110010011 : data = 16'b0101011010110001;
            15'b001010110010100 : data = 16'b0101011010011101;
            15'b001010110010101 : data = 16'b0101011010001010;
            15'b001010110010110 : data = 16'b0101011001110110;
            15'b001010110010111 : data = 16'b0101011001100011;
            15'b001010110011000 : data = 16'b0101011001001111;
            15'b001010110011001 : data = 16'b0101011000111100;
            15'b001010110011010 : data = 16'b0101011000101000;
            15'b001010110011011 : data = 16'b0101011000010101;
            15'b001010110011100 : data = 16'b0101011000000001;
            15'b001010110011101 : data = 16'b0101010111101110;
            15'b001010110011110 : data = 16'b0101010111011011;
            15'b001010110011111 : data = 16'b0101010111000111;
            15'b001010110100000 : data = 16'b0101010110110100;
            15'b001010110100001 : data = 16'b0101010110100000;
            15'b001010110100010 : data = 16'b0101010110001101;
            15'b001010110100011 : data = 16'b0101010101111001;
            15'b001010110100100 : data = 16'b0101010101100110;
            15'b001010110100101 : data = 16'b0101010101010011;
            15'b001010110100110 : data = 16'b0101010100111111;
            15'b001010110100111 : data = 16'b0101010100101100;
            15'b001010110101000 : data = 16'b0101010100011000;
            15'b001010110101001 : data = 16'b0101010100000101;
            15'b001010110101010 : data = 16'b0101010011110010;
            15'b001010110101011 : data = 16'b0101010011011110;
            15'b001010110101100 : data = 16'b0101010011001011;
            15'b001010110101101 : data = 16'b0101010010110111;
            15'b001010110101110 : data = 16'b0101010010100100;
            15'b001010110101111 : data = 16'b0101010010010001;
            15'b001010110110000 : data = 16'b0101010001111101;
            15'b001010110110001 : data = 16'b0101010001101010;
            15'b001010110110010 : data = 16'b0101010001010111;
            15'b001010110110011 : data = 16'b0101010001000011;
            15'b001010110110100 : data = 16'b0101010000110000;
            15'b001010110110101 : data = 16'b0101010000011101;
            15'b001010110110110 : data = 16'b0101010000001001;
            15'b001010110110111 : data = 16'b0101001111110110;
            15'b001010110111000 : data = 16'b0101001111100011;
            15'b001010110111001 : data = 16'b0101001111001111;
            15'b001010110111010 : data = 16'b0101001110111100;
            15'b001010110111011 : data = 16'b0101001110101001;
            15'b001010110111100 : data = 16'b0101001110010101;
            15'b001010110111101 : data = 16'b0101001110000010;
            15'b001010110111110 : data = 16'b0101001101101111;
            15'b001010110111111 : data = 16'b0101001101011011;
            15'b001010111000000 : data = 16'b0101001101001000;
            15'b001010111000001 : data = 16'b0101001100110101;
            15'b001010111000010 : data = 16'b0101001100100010;
            15'b001010111000011 : data = 16'b0101001100001110;
            15'b001010111000100 : data = 16'b0101001011111011;
            15'b001010111000101 : data = 16'b0101001011101000;
            15'b001010111000110 : data = 16'b0101001011010100;
            15'b001010111000111 : data = 16'b0101001011000001;
            15'b001010111001000 : data = 16'b0101001010101110;
            15'b001010111001001 : data = 16'b0101001010011011;
            15'b001010111001010 : data = 16'b0101001010000111;
            15'b001010111001011 : data = 16'b0101001001110100;
            15'b001010111001100 : data = 16'b0101001001100001;
            15'b001010111001101 : data = 16'b0101001001001110;
            15'b001010111001110 : data = 16'b0101001000111010;
            15'b001010111001111 : data = 16'b0101001000100111;
            15'b001010111010000 : data = 16'b0101001000010100;
            15'b001010111010001 : data = 16'b0101001000000001;
            15'b001010111010010 : data = 16'b0101000111101110;
            15'b001010111010011 : data = 16'b0101000111011010;
            15'b001010111010100 : data = 16'b0101000111000111;
            15'b001010111010101 : data = 16'b0101000110110100;
            15'b001010111010110 : data = 16'b0101000110100001;
            15'b001010111010111 : data = 16'b0101000110001110;
            15'b001010111011000 : data = 16'b0101000101111010;
            15'b001010111011001 : data = 16'b0101000101100111;
            15'b001010111011010 : data = 16'b0101000101010100;
            15'b001010111011011 : data = 16'b0101000101000001;
            15'b001010111011100 : data = 16'b0101000100101110;
            15'b001010111011101 : data = 16'b0101000100011011;
            15'b001010111011110 : data = 16'b0101000100000111;
            15'b001010111011111 : data = 16'b0101000011110100;
            15'b001010111100000 : data = 16'b0101000011100001;
            15'b001010111100001 : data = 16'b0101000011001110;
            15'b001010111100010 : data = 16'b0101000010111011;
            15'b001010111100011 : data = 16'b0101000010101000;
            15'b001010111100100 : data = 16'b0101000010010101;
            15'b001010111100101 : data = 16'b0101000010000010;
            15'b001010111100110 : data = 16'b0101000001101110;
            15'b001010111100111 : data = 16'b0101000001011011;
            15'b001010111101000 : data = 16'b0101000001001000;
            15'b001010111101001 : data = 16'b0101000000110101;
            15'b001010111101010 : data = 16'b0101000000100010;
            15'b001010111101011 : data = 16'b0101000000001111;
            15'b001010111101100 : data = 16'b0100111111111100;
            15'b001010111101101 : data = 16'b0100111111101001;
            15'b001010111101110 : data = 16'b0100111111010110;
            15'b001010111101111 : data = 16'b0100111111000011;
            15'b001010111110000 : data = 16'b0100111110101111;
            15'b001010111110001 : data = 16'b0100111110011100;
            15'b001010111110010 : data = 16'b0100111110001001;
            15'b001010111110011 : data = 16'b0100111101110110;
            15'b001010111110100 : data = 16'b0100111101100011;
            15'b001010111110101 : data = 16'b0100111101010000;
            15'b001010111110110 : data = 16'b0100111100111101;
            15'b001010111110111 : data = 16'b0100111100101010;
            15'b001010111111000 : data = 16'b0100111100010111;
            15'b001010111111001 : data = 16'b0100111100000100;
            15'b001010111111010 : data = 16'b0100111011110001;
            15'b001010111111011 : data = 16'b0100111011011110;
            15'b001010111111100 : data = 16'b0100111011001011;
            15'b001010111111101 : data = 16'b0100111010111000;
            15'b001010111111110 : data = 16'b0100111010100101;
            15'b001010111111111 : data = 16'b0100111010010010;
            15'b001011000000000 : data = 16'b0100111001111111;
            15'b001011000000001 : data = 16'b0100111001101100;
            15'b001011000000010 : data = 16'b0100111001011001;
            15'b001011000000011 : data = 16'b0100111001000110;
            15'b001011000000100 : data = 16'b0100111000110011;
            15'b001011000000101 : data = 16'b0100111000100000;
            15'b001011000000110 : data = 16'b0100111000001101;
            15'b001011000000111 : data = 16'b0100110111111010;
            15'b001011000001000 : data = 16'b0100110111100111;
            15'b001011000001001 : data = 16'b0100110111010100;
            15'b001011000001010 : data = 16'b0100110111000001;
            15'b001011000001011 : data = 16'b0100110110101111;
            15'b001011000001100 : data = 16'b0100110110011100;
            15'b001011000001101 : data = 16'b0100110110001001;
            15'b001011000001110 : data = 16'b0100110101110110;
            15'b001011000001111 : data = 16'b0100110101100011;
            15'b001011000010000 : data = 16'b0100110101010000;
            15'b001011000010001 : data = 16'b0100110100111101;
            15'b001011000010010 : data = 16'b0100110100101010;
            15'b001011000010011 : data = 16'b0100110100010111;
            15'b001011000010100 : data = 16'b0100110100000100;
            15'b001011000010101 : data = 16'b0100110011110001;
            15'b001011000010110 : data = 16'b0100110011011111;
            15'b001011000010111 : data = 16'b0100110011001100;
            15'b001011000011000 : data = 16'b0100110010111001;
            15'b001011000011001 : data = 16'b0100110010100110;
            15'b001011000011010 : data = 16'b0100110010010011;
            15'b001011000011011 : data = 16'b0100110010000000;
            15'b001011000011100 : data = 16'b0100110001101101;
            15'b001011000011101 : data = 16'b0100110001011011;
            15'b001011000011110 : data = 16'b0100110001001000;
            15'b001011000011111 : data = 16'b0100110000110101;
            15'b001011000100000 : data = 16'b0100110000100010;
            15'b001011000100001 : data = 16'b0100110000001111;
            15'b001011000100010 : data = 16'b0100101111111101;
            15'b001011000100011 : data = 16'b0100101111101010;
            15'b001011000100100 : data = 16'b0100101111010111;
            15'b001011000100101 : data = 16'b0100101111000100;
            15'b001011000100110 : data = 16'b0100101110110001;
            15'b001011000100111 : data = 16'b0100101110011111;
            15'b001011000101000 : data = 16'b0100101110001100;
            15'b001011000101001 : data = 16'b0100101101111001;
            15'b001011000101010 : data = 16'b0100101101100110;
            15'b001011000101011 : data = 16'b0100101101010011;
            15'b001011000101100 : data = 16'b0100101101000001;
            15'b001011000101101 : data = 16'b0100101100101110;
            15'b001011000101110 : data = 16'b0100101100011011;
            15'b001011000101111 : data = 16'b0100101100001000;
            15'b001011000110000 : data = 16'b0100101011110110;
            15'b001011000110001 : data = 16'b0100101011100011;
            15'b001011000110010 : data = 16'b0100101011010000;
            15'b001011000110011 : data = 16'b0100101010111101;
            15'b001011000110100 : data = 16'b0100101010101011;
            15'b001011000110101 : data = 16'b0100101010011000;
            15'b001011000110110 : data = 16'b0100101010000101;
            15'b001011000110111 : data = 16'b0100101001110011;
            15'b001011000111000 : data = 16'b0100101001100000;
            15'b001011000111001 : data = 16'b0100101001001101;
            15'b001011000111010 : data = 16'b0100101000111011;
            15'b001011000111011 : data = 16'b0100101000101000;
            15'b001011000111100 : data = 16'b0100101000010101;
            15'b001011000111101 : data = 16'b0100101000000011;
            15'b001011000111110 : data = 16'b0100100111110000;
            15'b001011000111111 : data = 16'b0100100111011101;
            15'b001011001000000 : data = 16'b0100100111001011;
            15'b001011001000001 : data = 16'b0100100110111000;
            15'b001011001000010 : data = 16'b0100100110100101;
            15'b001011001000011 : data = 16'b0100100110010011;
            15'b001011001000100 : data = 16'b0100100110000000;
            15'b001011001000101 : data = 16'b0100100101101101;
            15'b001011001000110 : data = 16'b0100100101011011;
            15'b001011001000111 : data = 16'b0100100101001000;
            15'b001011001001000 : data = 16'b0100100100110110;
            15'b001011001001001 : data = 16'b0100100100100011;
            15'b001011001001010 : data = 16'b0100100100010000;
            15'b001011001001011 : data = 16'b0100100011111110;
            15'b001011001001100 : data = 16'b0100100011101011;
            15'b001011001001101 : data = 16'b0100100011011001;
            15'b001011001001110 : data = 16'b0100100011000110;
            15'b001011001001111 : data = 16'b0100100010110011;
            15'b001011001010000 : data = 16'b0100100010100001;
            15'b001011001010001 : data = 16'b0100100010001110;
            15'b001011001010010 : data = 16'b0100100001111100;
            15'b001011001010011 : data = 16'b0100100001101001;
            15'b001011001010100 : data = 16'b0100100001010111;
            15'b001011001010101 : data = 16'b0100100001000100;
            15'b001011001010110 : data = 16'b0100100000110010;
            15'b001011001010111 : data = 16'b0100100000011111;
            15'b001011001011000 : data = 16'b0100100000001101;
            15'b001011001011001 : data = 16'b0100011111111010;
            15'b001011001011010 : data = 16'b0100011111101000;
            15'b001011001011011 : data = 16'b0100011111010101;
            15'b001011001011100 : data = 16'b0100011111000011;
            15'b001011001011101 : data = 16'b0100011110110000;
            15'b001011001011110 : data = 16'b0100011110011110;
            15'b001011001011111 : data = 16'b0100011110001011;
            15'b001011001100000 : data = 16'b0100011101111001;
            15'b001011001100001 : data = 16'b0100011101100110;
            15'b001011001100010 : data = 16'b0100011101010100;
            15'b001011001100011 : data = 16'b0100011101000001;
            15'b001011001100100 : data = 16'b0100011100101111;
            15'b001011001100101 : data = 16'b0100011100011100;
            15'b001011001100110 : data = 16'b0100011100001010;
            15'b001011001100111 : data = 16'b0100011011110111;
            15'b001011001101000 : data = 16'b0100011011100101;
            15'b001011001101001 : data = 16'b0100011011010011;
            15'b001011001101010 : data = 16'b0100011011000000;
            15'b001011001101011 : data = 16'b0100011010101110;
            15'b001011001101100 : data = 16'b0100011010011011;
            15'b001011001101101 : data = 16'b0100011010001001;
            15'b001011001101110 : data = 16'b0100011001110111;
            15'b001011001101111 : data = 16'b0100011001100100;
            15'b001011001110000 : data = 16'b0100011001010010;
            15'b001011001110001 : data = 16'b0100011000111111;
            15'b001011001110010 : data = 16'b0100011000101101;
            15'b001011001110011 : data = 16'b0100011000011011;
            15'b001011001110100 : data = 16'b0100011000001000;
            15'b001011001110101 : data = 16'b0100010111110110;
            15'b001011001110110 : data = 16'b0100010111100100;
            15'b001011001110111 : data = 16'b0100010111010001;
            15'b001011001111000 : data = 16'b0100010110111111;
            15'b001011001111001 : data = 16'b0100010110101101;
            15'b001011001111010 : data = 16'b0100010110011010;
            15'b001011001111011 : data = 16'b0100010110001000;
            15'b001011001111100 : data = 16'b0100010101110110;
            15'b001011001111101 : data = 16'b0100010101100011;
            15'b001011001111110 : data = 16'b0100010101010001;
            15'b001011001111111 : data = 16'b0100010100111111;
            15'b001011010000000 : data = 16'b0100010100101100;
            15'b001011010000001 : data = 16'b0100010100011010;
            15'b001011010000010 : data = 16'b0100010100001000;
            15'b001011010000011 : data = 16'b0100010011110110;
            15'b001011010000100 : data = 16'b0100010011100011;
            15'b001011010000101 : data = 16'b0100010011010001;
            15'b001011010000110 : data = 16'b0100010010111111;
            15'b001011010000111 : data = 16'b0100010010101101;
            15'b001011010001000 : data = 16'b0100010010011010;
            15'b001011010001001 : data = 16'b0100010010001000;
            15'b001011010001010 : data = 16'b0100010001110110;
            15'b001011010001011 : data = 16'b0100010001100100;
            15'b001011010001100 : data = 16'b0100010001010001;
            15'b001011010001101 : data = 16'b0100010000111111;
            15'b001011010001110 : data = 16'b0100010000101101;
            15'b001011010001111 : data = 16'b0100010000011011;
            15'b001011010010000 : data = 16'b0100010000001001;
            15'b001011010010001 : data = 16'b0100001111110110;
            15'b001011010010010 : data = 16'b0100001111100100;
            15'b001011010010011 : data = 16'b0100001111010010;
            15'b001011010010100 : data = 16'b0100001111000000;
            15'b001011010010101 : data = 16'b0100001110101110;
            15'b001011010010110 : data = 16'b0100001110011100;
            15'b001011010010111 : data = 16'b0100001110001001;
            15'b001011010011000 : data = 16'b0100001101110111;
            15'b001011010011001 : data = 16'b0100001101100101;
            15'b001011010011010 : data = 16'b0100001101010011;
            15'b001011010011011 : data = 16'b0100001101000001;
            15'b001011010011100 : data = 16'b0100001100101111;
            15'b001011010011101 : data = 16'b0100001100011101;
            15'b001011010011110 : data = 16'b0100001100001011;
            15'b001011010011111 : data = 16'b0100001011111001;
            15'b001011010100000 : data = 16'b0100001011100110;
            15'b001011010100001 : data = 16'b0100001011010100;
            15'b001011010100010 : data = 16'b0100001011000010;
            15'b001011010100011 : data = 16'b0100001010110000;
            15'b001011010100100 : data = 16'b0100001010011110;
            15'b001011010100101 : data = 16'b0100001010001100;
            15'b001011010100110 : data = 16'b0100001001111010;
            15'b001011010100111 : data = 16'b0100001001101000;
            15'b001011010101000 : data = 16'b0100001001010110;
            15'b001011010101001 : data = 16'b0100001001000100;
            15'b001011010101010 : data = 16'b0100001000110010;
            15'b001011010101011 : data = 16'b0100001000100000;
            15'b001011010101100 : data = 16'b0100001000001110;
            15'b001011010101101 : data = 16'b0100000111111100;
            15'b001011010101110 : data = 16'b0100000111101010;
            15'b001011010101111 : data = 16'b0100000111011000;
            15'b001011010110000 : data = 16'b0100000111000110;
            15'b001011010110001 : data = 16'b0100000110110100;
            15'b001011010110010 : data = 16'b0100000110100010;
            15'b001011010110011 : data = 16'b0100000110010000;
            15'b001011010110100 : data = 16'b0100000101111110;
            15'b001011010110101 : data = 16'b0100000101101100;
            15'b001011010110110 : data = 16'b0100000101011010;
            15'b001011010110111 : data = 16'b0100000101001000;
            15'b001011010111000 : data = 16'b0100000100110110;
            15'b001011010111001 : data = 16'b0100000100100100;
            15'b001011010111010 : data = 16'b0100000100010010;
            15'b001011010111011 : data = 16'b0100000100000000;
            15'b001011010111100 : data = 16'b0100000011101110;
            15'b001011010111101 : data = 16'b0100000011011100;
            15'b001011010111110 : data = 16'b0100000011001010;
            15'b001011010111111 : data = 16'b0100000010111001;
            15'b001011011000000 : data = 16'b0100000010100111;
            15'b001011011000001 : data = 16'b0100000010010101;
            15'b001011011000010 : data = 16'b0100000010000011;
            15'b001011011000011 : data = 16'b0100000001110001;
            15'b001011011000100 : data = 16'b0100000001011111;
            15'b001011011000101 : data = 16'b0100000001001101;
            15'b001011011000110 : data = 16'b0100000000111011;
            15'b001011011000111 : data = 16'b0100000000101010;
            15'b001011011001000 : data = 16'b0100000000011000;
            15'b001011011001001 : data = 16'b0100000000000110;
            15'b001011011001010 : data = 16'b0011111111110100;
            15'b001011011001011 : data = 16'b0011111111100010;
            15'b001011011001100 : data = 16'b0011111111010000;
            15'b001011011001101 : data = 16'b0011111110111111;
            15'b001011011001110 : data = 16'b0011111110101101;
            15'b001011011001111 : data = 16'b0011111110011011;
            15'b001011011010000 : data = 16'b0011111110001001;
            15'b001011011010001 : data = 16'b0011111101110111;
            15'b001011011010010 : data = 16'b0011111101100110;
            15'b001011011010011 : data = 16'b0011111101010100;
            15'b001011011010100 : data = 16'b0011111101000010;
            15'b001011011010101 : data = 16'b0011111100110000;
            15'b001011011010110 : data = 16'b0011111100011111;
            15'b001011011010111 : data = 16'b0011111100001101;
            15'b001011011011000 : data = 16'b0011111011111011;
            15'b001011011011001 : data = 16'b0011111011101001;
            15'b001011011011010 : data = 16'b0011111011011000;
            15'b001011011011011 : data = 16'b0011111011000110;
            15'b001011011011100 : data = 16'b0011111010110100;
            15'b001011011011101 : data = 16'b0011111010100011;
            15'b001011011011110 : data = 16'b0011111010010001;
            15'b001011011011111 : data = 16'b0011111001111111;
            15'b001011011100000 : data = 16'b0011111001101110;
            15'b001011011100001 : data = 16'b0011111001011100;
            15'b001011011100010 : data = 16'b0011111001001010;
            15'b001011011100011 : data = 16'b0011111000111001;
            15'b001011011100100 : data = 16'b0011111000100111;
            15'b001011011100101 : data = 16'b0011111000010101;
            15'b001011011100110 : data = 16'b0011111000000100;
            15'b001011011100111 : data = 16'b0011110111110010;
            15'b001011011101000 : data = 16'b0011110111100000;
            15'b001011011101001 : data = 16'b0011110111001111;
            15'b001011011101010 : data = 16'b0011110110111101;
            15'b001011011101011 : data = 16'b0011110110101011;
            15'b001011011101100 : data = 16'b0011110110011010;
            15'b001011011101101 : data = 16'b0011110110001000;
            15'b001011011101110 : data = 16'b0011110101110111;
            15'b001011011101111 : data = 16'b0011110101100101;
            15'b001011011110000 : data = 16'b0011110101010011;
            15'b001011011110001 : data = 16'b0011110101000010;
            15'b001011011110010 : data = 16'b0011110100110000;
            15'b001011011110011 : data = 16'b0011110100011111;
            15'b001011011110100 : data = 16'b0011110100001101;
            15'b001011011110101 : data = 16'b0011110011111100;
            15'b001011011110110 : data = 16'b0011110011101010;
            15'b001011011110111 : data = 16'b0011110011011001;
            15'b001011011111000 : data = 16'b0011110011000111;
            15'b001011011111001 : data = 16'b0011110010110110;
            15'b001011011111010 : data = 16'b0011110010100100;
            15'b001011011111011 : data = 16'b0011110010010011;
            15'b001011011111100 : data = 16'b0011110010000001;
            15'b001011011111101 : data = 16'b0011110001110000;
            15'b001011011111110 : data = 16'b0011110001011110;
            15'b001011011111111 : data = 16'b0011110001001101;
            15'b001011100000000 : data = 16'b0011110000111011;
            15'b001011100000001 : data = 16'b0011110000101010;
            15'b001011100000010 : data = 16'b0011110000011000;
            15'b001011100000011 : data = 16'b0011110000000111;
            15'b001011100000100 : data = 16'b0011101111110101;
            15'b001011100000101 : data = 16'b0011101111100100;
            15'b001011100000110 : data = 16'b0011101111010010;
            15'b001011100000111 : data = 16'b0011101111000001;
            15'b001011100001000 : data = 16'b0011101110110000;
            15'b001011100001001 : data = 16'b0011101110011110;
            15'b001011100001010 : data = 16'b0011101110001101;
            15'b001011100001011 : data = 16'b0011101101111011;
            15'b001011100001100 : data = 16'b0011101101101010;
            15'b001011100001101 : data = 16'b0011101101011001;
            15'b001011100001110 : data = 16'b0011101101000111;
            15'b001011100001111 : data = 16'b0011101100110110;
            15'b001011100010000 : data = 16'b0011101100100101;
            15'b001011100010001 : data = 16'b0011101100010011;
            15'b001011100010010 : data = 16'b0011101100000010;
            15'b001011100010011 : data = 16'b0011101011110001;
            15'b001011100010100 : data = 16'b0011101011011111;
            15'b001011100010101 : data = 16'b0011101011001110;
            15'b001011100010110 : data = 16'b0011101010111101;
            15'b001011100010111 : data = 16'b0011101010101011;
            15'b001011100011000 : data = 16'b0011101010011010;
            15'b001011100011001 : data = 16'b0011101010001001;
            15'b001011100011010 : data = 16'b0011101001110111;
            15'b001011100011011 : data = 16'b0011101001100110;
            15'b001011100011100 : data = 16'b0011101001010101;
            15'b001011100011101 : data = 16'b0011101001000100;
            15'b001011100011110 : data = 16'b0011101000110010;
            15'b001011100011111 : data = 16'b0011101000100001;
            15'b001011100100000 : data = 16'b0011101000010000;
            15'b001011100100001 : data = 16'b0011100111111111;
            15'b001011100100010 : data = 16'b0011100111101101;
            15'b001011100100011 : data = 16'b0011100111011100;
            15'b001011100100100 : data = 16'b0011100111001011;
            15'b001011100100101 : data = 16'b0011100110111010;
            15'b001011100100110 : data = 16'b0011100110101000;
            15'b001011100100111 : data = 16'b0011100110010111;
            15'b001011100101000 : data = 16'b0011100110000110;
            15'b001011100101001 : data = 16'b0011100101110101;
            15'b001011100101010 : data = 16'b0011100101100100;
            15'b001011100101011 : data = 16'b0011100101010011;
            15'b001011100101100 : data = 16'b0011100101000001;
            15'b001011100101101 : data = 16'b0011100100110000;
            15'b001011100101110 : data = 16'b0011100100011111;
            15'b001011100101111 : data = 16'b0011100100001110;
            15'b001011100110000 : data = 16'b0011100011111101;
            15'b001011100110001 : data = 16'b0011100011101100;
            15'b001011100110010 : data = 16'b0011100011011011;
            15'b001011100110011 : data = 16'b0011100011001001;
            15'b001011100110100 : data = 16'b0011100010111000;
            15'b001011100110101 : data = 16'b0011100010100111;
            15'b001011100110110 : data = 16'b0011100010010110;
            15'b001011100110111 : data = 16'b0011100010000101;
            15'b001011100111000 : data = 16'b0011100001110100;
            15'b001011100111001 : data = 16'b0011100001100011;
            15'b001011100111010 : data = 16'b0011100001010010;
            15'b001011100111011 : data = 16'b0011100001000001;
            15'b001011100111100 : data = 16'b0011100000110000;
            15'b001011100111101 : data = 16'b0011100000011111;
            15'b001011100111110 : data = 16'b0011100000001110;
            15'b001011100111111 : data = 16'b0011011111111101;
            15'b001011101000000 : data = 16'b0011011111101100;
            15'b001011101000001 : data = 16'b0011011111011011;
            15'b001011101000010 : data = 16'b0011011111001010;
            15'b001011101000011 : data = 16'b0011011110111001;
            15'b001011101000100 : data = 16'b0011011110101000;
            15'b001011101000101 : data = 16'b0011011110010111;
            15'b001011101000110 : data = 16'b0011011110000110;
            15'b001011101000111 : data = 16'b0011011101110101;
            15'b001011101001000 : data = 16'b0011011101100100;
            15'b001011101001001 : data = 16'b0011011101010011;
            15'b001011101001010 : data = 16'b0011011101000010;
            15'b001011101001011 : data = 16'b0011011100110001;
            15'b001011101001100 : data = 16'b0011011100100000;
            15'b001011101001101 : data = 16'b0011011100001111;
            15'b001011101001110 : data = 16'b0011011011111110;
            15'b001011101001111 : data = 16'b0011011011101101;
            15'b001011101010000 : data = 16'b0011011011011100;
            15'b001011101010001 : data = 16'b0011011011001100;
            15'b001011101010010 : data = 16'b0011011010111011;
            15'b001011101010011 : data = 16'b0011011010101010;
            15'b001011101010100 : data = 16'b0011011010011001;
            15'b001011101010101 : data = 16'b0011011010001000;
            15'b001011101010110 : data = 16'b0011011001110111;
            15'b001011101010111 : data = 16'b0011011001100110;
            15'b001011101011000 : data = 16'b0011011001010101;
            15'b001011101011001 : data = 16'b0011011001000101;
            15'b001011101011010 : data = 16'b0011011000110100;
            15'b001011101011011 : data = 16'b0011011000100011;
            15'b001011101011100 : data = 16'b0011011000010010;
            15'b001011101011101 : data = 16'b0011011000000001;
            15'b001011101011110 : data = 16'b0011010111110001;
            15'b001011101011111 : data = 16'b0011010111100000;
            15'b001011101100000 : data = 16'b0011010111001111;
            15'b001011101100001 : data = 16'b0011010110111110;
            15'b001011101100010 : data = 16'b0011010110101101;
            15'b001011101100011 : data = 16'b0011010110011101;
            15'b001011101100100 : data = 16'b0011010110001100;
            15'b001011101100101 : data = 16'b0011010101111011;
            15'b001011101100110 : data = 16'b0011010101101010;
            15'b001011101100111 : data = 16'b0011010101011010;
            15'b001011101101000 : data = 16'b0011010101001001;
            15'b001011101101001 : data = 16'b0011010100111000;
            15'b001011101101010 : data = 16'b0011010100101000;
            15'b001011101101011 : data = 16'b0011010100010111;
            15'b001011101101100 : data = 16'b0011010100000110;
            15'b001011101101101 : data = 16'b0011010011110110;
            15'b001011101101110 : data = 16'b0011010011100101;
            15'b001011101101111 : data = 16'b0011010011010100;
            15'b001011101110000 : data = 16'b0011010011000100;
            15'b001011101110001 : data = 16'b0011010010110011;
            15'b001011101110010 : data = 16'b0011010010100010;
            15'b001011101110011 : data = 16'b0011010010010010;
            15'b001011101110100 : data = 16'b0011010010000001;
            15'b001011101110101 : data = 16'b0011010001110000;
            15'b001011101110110 : data = 16'b0011010001100000;
            15'b001011101110111 : data = 16'b0011010001001111;
            15'b001011101111000 : data = 16'b0011010000111111;
            15'b001011101111001 : data = 16'b0011010000101110;
            15'b001011101111010 : data = 16'b0011010000011101;
            15'b001011101111011 : data = 16'b0011010000001101;
            15'b001011101111100 : data = 16'b0011001111111100;
            15'b001011101111101 : data = 16'b0011001111101100;
            15'b001011101111110 : data = 16'b0011001111011011;
            15'b001011101111111 : data = 16'b0011001111001011;
            15'b001011110000000 : data = 16'b0011001110111010;
            15'b001011110000001 : data = 16'b0011001110101001;
            15'b001011110000010 : data = 16'b0011001110011001;
            15'b001011110000011 : data = 16'b0011001110001000;
            15'b001011110000100 : data = 16'b0011001101111000;
            15'b001011110000101 : data = 16'b0011001101100111;
            15'b001011110000110 : data = 16'b0011001101010111;
            15'b001011110000111 : data = 16'b0011001101000110;
            15'b001011110001000 : data = 16'b0011001100110110;
            15'b001011110001001 : data = 16'b0011001100100110;
            15'b001011110001010 : data = 16'b0011001100010101;
            15'b001011110001011 : data = 16'b0011001100000101;
            15'b001011110001100 : data = 16'b0011001011110100;
            15'b001011110001101 : data = 16'b0011001011100100;
            15'b001011110001110 : data = 16'b0011001011010011;
            15'b001011110001111 : data = 16'b0011001011000011;
            15'b001011110010000 : data = 16'b0011001010110010;
            15'b001011110010001 : data = 16'b0011001010100010;
            15'b001011110010010 : data = 16'b0011001010010010;
            15'b001011110010011 : data = 16'b0011001010000001;
            15'b001011110010100 : data = 16'b0011001001110001;
            15'b001011110010101 : data = 16'b0011001001100001;
            15'b001011110010110 : data = 16'b0011001001010000;
            15'b001011110010111 : data = 16'b0011001001000000;
            15'b001011110011000 : data = 16'b0011001000101111;
            15'b001011110011001 : data = 16'b0011001000011111;
            15'b001011110011010 : data = 16'b0011001000001111;
            15'b001011110011011 : data = 16'b0011000111111110;
            15'b001011110011100 : data = 16'b0011000111101110;
            15'b001011110011101 : data = 16'b0011000111011110;
            15'b001011110011110 : data = 16'b0011000111001110;
            15'b001011110011111 : data = 16'b0011000110111101;
            15'b001011110100000 : data = 16'b0011000110101101;
            15'b001011110100001 : data = 16'b0011000110011101;
            15'b001011110100010 : data = 16'b0011000110001100;
            15'b001011110100011 : data = 16'b0011000101111100;
            15'b001011110100100 : data = 16'b0011000101101100;
            15'b001011110100101 : data = 16'b0011000101011100;
            15'b001011110100110 : data = 16'b0011000101001011;
            15'b001011110100111 : data = 16'b0011000100111011;
            15'b001011110101000 : data = 16'b0011000100101011;
            15'b001011110101001 : data = 16'b0011000100011011;
            15'b001011110101010 : data = 16'b0011000100001010;
            15'b001011110101011 : data = 16'b0011000011111010;
            15'b001011110101100 : data = 16'b0011000011101010;
            15'b001011110101101 : data = 16'b0011000011011010;
            15'b001011110101110 : data = 16'b0011000011001010;
            15'b001011110101111 : data = 16'b0011000010111010;
            15'b001011110110000 : data = 16'b0011000010101001;
            15'b001011110110001 : data = 16'b0011000010011001;
            15'b001011110110010 : data = 16'b0011000010001001;
            15'b001011110110011 : data = 16'b0011000001111001;
            15'b001011110110100 : data = 16'b0011000001101001;
            15'b001011110110101 : data = 16'b0011000001011001;
            15'b001011110110110 : data = 16'b0011000001001001;
            15'b001011110110111 : data = 16'b0011000000111001;
            15'b001011110111000 : data = 16'b0011000000101000;
            15'b001011110111001 : data = 16'b0011000000011000;
            15'b001011110111010 : data = 16'b0011000000001000;
            15'b001011110111011 : data = 16'b0010111111111000;
            15'b001011110111100 : data = 16'b0010111111101000;
            15'b001011110111101 : data = 16'b0010111111011000;
            15'b001011110111110 : data = 16'b0010111111001000;
            15'b001011110111111 : data = 16'b0010111110111000;
            15'b001011111000000 : data = 16'b0010111110101000;
            15'b001011111000001 : data = 16'b0010111110011000;
            15'b001011111000010 : data = 16'b0010111110001000;
            15'b001011111000011 : data = 16'b0010111101111000;
            15'b001011111000100 : data = 16'b0010111101101000;
            15'b001011111000101 : data = 16'b0010111101011000;
            15'b001011111000110 : data = 16'b0010111101001000;
            15'b001011111000111 : data = 16'b0010111100111000;
            15'b001011111001000 : data = 16'b0010111100101000;
            15'b001011111001001 : data = 16'b0010111100011000;
            15'b001011111001010 : data = 16'b0010111100001000;
            15'b001011111001011 : data = 16'b0010111011111000;
            15'b001011111001100 : data = 16'b0010111011101000;
            15'b001011111001101 : data = 16'b0010111011011000;
            15'b001011111001110 : data = 16'b0010111011001000;
            15'b001011111001111 : data = 16'b0010111010111000;
            15'b001011111010000 : data = 16'b0010111010101001;
            15'b001011111010001 : data = 16'b0010111010011001;
            15'b001011111010010 : data = 16'b0010111010001001;
            15'b001011111010011 : data = 16'b0010111001111001;
            15'b001011111010100 : data = 16'b0010111001101001;
            15'b001011111010101 : data = 16'b0010111001011001;
            15'b001011111010110 : data = 16'b0010111001001001;
            15'b001011111010111 : data = 16'b0010111000111001;
            15'b001011111011000 : data = 16'b0010111000101010;
            15'b001011111011001 : data = 16'b0010111000011010;
            15'b001011111011010 : data = 16'b0010111000001010;
            15'b001011111011011 : data = 16'b0010110111111010;
            15'b001011111011100 : data = 16'b0010110111101010;
            15'b001011111011101 : data = 16'b0010110111011011;
            15'b001011111011110 : data = 16'b0010110111001011;
            15'b001011111011111 : data = 16'b0010110110111011;
            15'b001011111100000 : data = 16'b0010110110101011;
            15'b001011111100001 : data = 16'b0010110110011100;
            15'b001011111100010 : data = 16'b0010110110001100;
            15'b001011111100011 : data = 16'b0010110101111100;
            15'b001011111100100 : data = 16'b0010110101101100;
            15'b001011111100101 : data = 16'b0010110101011101;
            15'b001011111100110 : data = 16'b0010110101001101;
            15'b001011111100111 : data = 16'b0010110100111101;
            15'b001011111101000 : data = 16'b0010110100101101;
            15'b001011111101001 : data = 16'b0010110100011110;
            15'b001011111101010 : data = 16'b0010110100001110;
            15'b001011111101011 : data = 16'b0010110011111110;
            15'b001011111101100 : data = 16'b0010110011101111;
            15'b001011111101101 : data = 16'b0010110011011111;
            15'b001011111101110 : data = 16'b0010110011001111;
            15'b001011111101111 : data = 16'b0010110011000000;
            15'b001011111110000 : data = 16'b0010110010110000;
            15'b001011111110001 : data = 16'b0010110010100000;
            15'b001011111110010 : data = 16'b0010110010010001;
            15'b001011111110011 : data = 16'b0010110010000001;
            15'b001011111110100 : data = 16'b0010110001110010;
            15'b001011111110101 : data = 16'b0010110001100010;
            15'b001011111110110 : data = 16'b0010110001010010;
            15'b001011111110111 : data = 16'b0010110001000011;
            15'b001011111111000 : data = 16'b0010110000110011;
            15'b001011111111001 : data = 16'b0010110000100100;
            15'b001011111111010 : data = 16'b0010110000010100;
            15'b001011111111011 : data = 16'b0010110000000101;
            15'b001011111111100 : data = 16'b0010101111110101;
            15'b001011111111101 : data = 16'b0010101111100110;
            15'b001011111111110 : data = 16'b0010101111010110;
            15'b001011111111111 : data = 16'b0010101111000111;
            15'b001100000000000 : data = 16'b0010101110110111;
            15'b001100000000001 : data = 16'b0010101110101000;
            15'b001100000000010 : data = 16'b0010101110011000;
            15'b001100000000011 : data = 16'b0010101110001001;
            15'b001100000000100 : data = 16'b0010101101111001;
            15'b001100000000101 : data = 16'b0010101101101010;
            15'b001100000000110 : data = 16'b0010101101011010;
            15'b001100000000111 : data = 16'b0010101101001011;
            15'b001100000001000 : data = 16'b0010101100111011;
            15'b001100000001001 : data = 16'b0010101100101100;
            15'b001100000001010 : data = 16'b0010101100011101;
            15'b001100000001011 : data = 16'b0010101100001101;
            15'b001100000001100 : data = 16'b0010101011111110;
            15'b001100000001101 : data = 16'b0010101011101110;
            15'b001100000001110 : data = 16'b0010101011011111;
            15'b001100000001111 : data = 16'b0010101011010000;
            15'b001100000010000 : data = 16'b0010101011000000;
            15'b001100000010001 : data = 16'b0010101010110001;
            15'b001100000010010 : data = 16'b0010101010100010;
            15'b001100000010011 : data = 16'b0010101010010010;
            15'b001100000010100 : data = 16'b0010101010000011;
            15'b001100000010101 : data = 16'b0010101001110100;
            15'b001100000010110 : data = 16'b0010101001100100;
            15'b001100000010111 : data = 16'b0010101001010101;
            15'b001100000011000 : data = 16'b0010101001000110;
            15'b001100000011001 : data = 16'b0010101000110110;
            15'b001100000011010 : data = 16'b0010101000100111;
            15'b001100000011011 : data = 16'b0010101000011000;
            15'b001100000011100 : data = 16'b0010101000001001;
            15'b001100000011101 : data = 16'b0010100111111001;
            15'b001100000011110 : data = 16'b0010100111101010;
            15'b001100000011111 : data = 16'b0010100111011011;
            15'b001100000100000 : data = 16'b0010100111001100;
            15'b001100000100001 : data = 16'b0010100110111100;
            15'b001100000100010 : data = 16'b0010100110101101;
            15'b001100000100011 : data = 16'b0010100110011110;
            15'b001100000100100 : data = 16'b0010100110001111;
            15'b001100000100101 : data = 16'b0010100110000000;
            15'b001100000100110 : data = 16'b0010100101110001;
            15'b001100000100111 : data = 16'b0010100101100001;
            15'b001100000101000 : data = 16'b0010100101010010;
            15'b001100000101001 : data = 16'b0010100101000011;
            15'b001100000101010 : data = 16'b0010100100110100;
            15'b001100000101011 : data = 16'b0010100100100101;
            15'b001100000101100 : data = 16'b0010100100010110;
            15'b001100000101101 : data = 16'b0010100100000111;
            15'b001100000101110 : data = 16'b0010100011110111;
            15'b001100000101111 : data = 16'b0010100011101000;
            15'b001100000110000 : data = 16'b0010100011011001;
            15'b001100000110001 : data = 16'b0010100011001010;
            15'b001100000110010 : data = 16'b0010100010111011;
            15'b001100000110011 : data = 16'b0010100010101100;
            15'b001100000110100 : data = 16'b0010100010011101;
            15'b001100000110101 : data = 16'b0010100010001110;
            15'b001100000110110 : data = 16'b0010100001111111;
            15'b001100000110111 : data = 16'b0010100001110000;
            15'b001100000111000 : data = 16'b0010100001100001;
            15'b001100000111001 : data = 16'b0010100001010010;
            15'b001100000111010 : data = 16'b0010100001000011;
            15'b001100000111011 : data = 16'b0010100000110100;
            15'b001100000111100 : data = 16'b0010100000100101;
            15'b001100000111101 : data = 16'b0010100000010110;
            15'b001100000111110 : data = 16'b0010100000000111;
            15'b001100000111111 : data = 16'b0010011111111000;
            15'b001100001000000 : data = 16'b0010011111101001;
            15'b001100001000001 : data = 16'b0010011111011010;
            15'b001100001000010 : data = 16'b0010011111001011;
            15'b001100001000011 : data = 16'b0010011110111100;
            15'b001100001000100 : data = 16'b0010011110101101;
            15'b001100001000101 : data = 16'b0010011110011111;
            15'b001100001000110 : data = 16'b0010011110010000;
            15'b001100001000111 : data = 16'b0010011110000001;
            15'b001100001001000 : data = 16'b0010011101110010;
            15'b001100001001001 : data = 16'b0010011101100011;
            15'b001100001001010 : data = 16'b0010011101010100;
            15'b001100001001011 : data = 16'b0010011101000101;
            15'b001100001001100 : data = 16'b0010011100110111;
            15'b001100001001101 : data = 16'b0010011100101000;
            15'b001100001001110 : data = 16'b0010011100011001;
            15'b001100001001111 : data = 16'b0010011100001010;
            15'b001100001010000 : data = 16'b0010011011111011;
            15'b001100001010001 : data = 16'b0010011011101101;
            15'b001100001010010 : data = 16'b0010011011011110;
            15'b001100001010011 : data = 16'b0010011011001111;
            15'b001100001010100 : data = 16'b0010011011000000;
            15'b001100001010101 : data = 16'b0010011010110001;
            15'b001100001010110 : data = 16'b0010011010100011;
            15'b001100001010111 : data = 16'b0010011010010100;
            15'b001100001011000 : data = 16'b0010011010000101;
            15'b001100001011001 : data = 16'b0010011001110111;
            15'b001100001011010 : data = 16'b0010011001101000;
            15'b001100001011011 : data = 16'b0010011001011001;
            15'b001100001011100 : data = 16'b0010011001001010;
            15'b001100001011101 : data = 16'b0010011000111100;
            15'b001100001011110 : data = 16'b0010011000101101;
            15'b001100001011111 : data = 16'b0010011000011110;
            15'b001100001100000 : data = 16'b0010011000010000;
            15'b001100001100001 : data = 16'b0010011000000001;
            15'b001100001100010 : data = 16'b0010010111110010;
            15'b001100001100011 : data = 16'b0010010111100100;
            15'b001100001100100 : data = 16'b0010010111010101;
            15'b001100001100101 : data = 16'b0010010111000111;
            15'b001100001100110 : data = 16'b0010010110111000;
            15'b001100001100111 : data = 16'b0010010110101001;
            15'b001100001101000 : data = 16'b0010010110011011;
            15'b001100001101001 : data = 16'b0010010110001100;
            15'b001100001101010 : data = 16'b0010010101111110;
            15'b001100001101011 : data = 16'b0010010101101111;
            15'b001100001101100 : data = 16'b0010010101100001;
            15'b001100001101101 : data = 16'b0010010101010010;
            15'b001100001101110 : data = 16'b0010010101000100;
            15'b001100001101111 : data = 16'b0010010100110101;
            15'b001100001110000 : data = 16'b0010010100100111;
            15'b001100001110001 : data = 16'b0010010100011000;
            15'b001100001110010 : data = 16'b0010010100001010;
            15'b001100001110011 : data = 16'b0010010011111011;
            15'b001100001110100 : data = 16'b0010010011101101;
            15'b001100001110101 : data = 16'b0010010011011110;
            15'b001100001110110 : data = 16'b0010010011010000;
            15'b001100001110111 : data = 16'b0010010011000001;
            15'b001100001111000 : data = 16'b0010010010110011;
            15'b001100001111001 : data = 16'b0010010010100100;
            15'b001100001111010 : data = 16'b0010010010010110;
            15'b001100001111011 : data = 16'b0010010010001000;
            15'b001100001111100 : data = 16'b0010010001111001;
            15'b001100001111101 : data = 16'b0010010001101011;
            15'b001100001111110 : data = 16'b0010010001011100;
            15'b001100001111111 : data = 16'b0010010001001110;
            15'b001100010000000 : data = 16'b0010010001000000;
            15'b001100010000001 : data = 16'b0010010000110001;
            15'b001100010000010 : data = 16'b0010010000100011;
            15'b001100010000011 : data = 16'b0010010000010101;
            15'b001100010000100 : data = 16'b0010010000000110;
            15'b001100010000101 : data = 16'b0010001111111000;
            15'b001100010000110 : data = 16'b0010001111101010;
            15'b001100010000111 : data = 16'b0010001111011011;
            15'b001100010001000 : data = 16'b0010001111001101;
            15'b001100010001001 : data = 16'b0010001110111111;
            15'b001100010001010 : data = 16'b0010001110110001;
            15'b001100010001011 : data = 16'b0010001110100010;
            15'b001100010001100 : data = 16'b0010001110010100;
            15'b001100010001101 : data = 16'b0010001110000110;
            15'b001100010001110 : data = 16'b0010001101111000;
            15'b001100010001111 : data = 16'b0010001101101001;
            15'b001100010010000 : data = 16'b0010001101011011;
            15'b001100010010001 : data = 16'b0010001101001101;
            15'b001100010010010 : data = 16'b0010001100111111;
            15'b001100010010011 : data = 16'b0010001100110001;
            15'b001100010010100 : data = 16'b0010001100100010;
            15'b001100010010101 : data = 16'b0010001100010100;
            15'b001100010010110 : data = 16'b0010001100000110;
            15'b001100010010111 : data = 16'b0010001011111000;
            15'b001100010011000 : data = 16'b0010001011101010;
            15'b001100010011001 : data = 16'b0010001011011100;
            15'b001100010011010 : data = 16'b0010001011001110;
            15'b001100010011011 : data = 16'b0010001010111111;
            15'b001100010011100 : data = 16'b0010001010110001;
            15'b001100010011101 : data = 16'b0010001010100011;
            15'b001100010011110 : data = 16'b0010001010010101;
            15'b001100010011111 : data = 16'b0010001010000111;
            15'b001100010100000 : data = 16'b0010001001111001;
            15'b001100010100001 : data = 16'b0010001001101011;
            15'b001100010100010 : data = 16'b0010001001011101;
            15'b001100010100011 : data = 16'b0010001001001111;
            15'b001100010100100 : data = 16'b0010001001000001;
            15'b001100010100101 : data = 16'b0010001000110011;
            15'b001100010100110 : data = 16'b0010001000100101;
            15'b001100010100111 : data = 16'b0010001000010111;
            15'b001100010101000 : data = 16'b0010001000001001;
            15'b001100010101001 : data = 16'b0010000111111011;
            15'b001100010101010 : data = 16'b0010000111101101;
            15'b001100010101011 : data = 16'b0010000111011111;
            15'b001100010101100 : data = 16'b0010000111010001;
            15'b001100010101101 : data = 16'b0010000111000011;
            15'b001100010101110 : data = 16'b0010000110110101;
            15'b001100010101111 : data = 16'b0010000110100111;
            15'b001100010110000 : data = 16'b0010000110011001;
            15'b001100010110001 : data = 16'b0010000110001100;
            15'b001100010110010 : data = 16'b0010000101111110;
            15'b001100010110011 : data = 16'b0010000101110000;
            15'b001100010110100 : data = 16'b0010000101100010;
            15'b001100010110101 : data = 16'b0010000101010100;
            15'b001100010110110 : data = 16'b0010000101000110;
            15'b001100010110111 : data = 16'b0010000100111000;
            15'b001100010111000 : data = 16'b0010000100101010;
            15'b001100010111001 : data = 16'b0010000100011101;
            15'b001100010111010 : data = 16'b0010000100001111;
            15'b001100010111011 : data = 16'b0010000100000001;
            15'b001100010111100 : data = 16'b0010000011110011;
            15'b001100010111101 : data = 16'b0010000011100101;
            15'b001100010111110 : data = 16'b0010000011011000;
            15'b001100010111111 : data = 16'b0010000011001010;
            15'b001100011000000 : data = 16'b0010000010111100;
            15'b001100011000001 : data = 16'b0010000010101110;
            15'b001100011000010 : data = 16'b0010000010100001;
            15'b001100011000011 : data = 16'b0010000010010011;
            15'b001100011000100 : data = 16'b0010000010000101;
            15'b001100011000101 : data = 16'b0010000001111000;
            15'b001100011000110 : data = 16'b0010000001101010;
            15'b001100011000111 : data = 16'b0010000001011100;
            15'b001100011001000 : data = 16'b0010000001001110;
            15'b001100011001001 : data = 16'b0010000001000001;
            15'b001100011001010 : data = 16'b0010000000110011;
            15'b001100011001011 : data = 16'b0010000000100101;
            15'b001100011001100 : data = 16'b0010000000011000;
            15'b001100011001101 : data = 16'b0010000000001010;
            15'b001100011001110 : data = 16'b0001111111111101;
            15'b001100011001111 : data = 16'b0001111111101111;
            15'b001100011010000 : data = 16'b0001111111100001;
            15'b001100011010001 : data = 16'b0001111111010100;
            15'b001100011010010 : data = 16'b0001111111000110;
            15'b001100011010011 : data = 16'b0001111110111001;
            15'b001100011010100 : data = 16'b0001111110101011;
            15'b001100011010101 : data = 16'b0001111110011110;
            15'b001100011010110 : data = 16'b0001111110010000;
            15'b001100011010111 : data = 16'b0001111110000010;
            15'b001100011011000 : data = 16'b0001111101110101;
            15'b001100011011001 : data = 16'b0001111101100111;
            15'b001100011011010 : data = 16'b0001111101011010;
            15'b001100011011011 : data = 16'b0001111101001100;
            15'b001100011011100 : data = 16'b0001111100111111;
            15'b001100011011101 : data = 16'b0001111100110001;
            15'b001100011011110 : data = 16'b0001111100100100;
            15'b001100011011111 : data = 16'b0001111100010111;
            15'b001100011100000 : data = 16'b0001111100001001;
            15'b001100011100001 : data = 16'b0001111011111100;
            15'b001100011100010 : data = 16'b0001111011101110;
            15'b001100011100011 : data = 16'b0001111011100001;
            15'b001100011100100 : data = 16'b0001111011010011;
            15'b001100011100101 : data = 16'b0001111011000110;
            15'b001100011100110 : data = 16'b0001111010111001;
            15'b001100011100111 : data = 16'b0001111010101011;
            15'b001100011101000 : data = 16'b0001111010011110;
            15'b001100011101001 : data = 16'b0001111010010001;
            15'b001100011101010 : data = 16'b0001111010000011;
            15'b001100011101011 : data = 16'b0001111001110110;
            15'b001100011101100 : data = 16'b0001111001101001;
            15'b001100011101101 : data = 16'b0001111001011011;
            15'b001100011101110 : data = 16'b0001111001001110;
            15'b001100011101111 : data = 16'b0001111001000001;
            15'b001100011110000 : data = 16'b0001111000110011;
            15'b001100011110001 : data = 16'b0001111000100110;
            15'b001100011110010 : data = 16'b0001111000011001;
            15'b001100011110011 : data = 16'b0001111000001100;
            15'b001100011110100 : data = 16'b0001110111111110;
            15'b001100011110101 : data = 16'b0001110111110001;
            15'b001100011110110 : data = 16'b0001110111100100;
            15'b001100011110111 : data = 16'b0001110111010111;
            15'b001100011111000 : data = 16'b0001110111001001;
            15'b001100011111001 : data = 16'b0001110110111100;
            15'b001100011111010 : data = 16'b0001110110101111;
            15'b001100011111011 : data = 16'b0001110110100010;
            15'b001100011111100 : data = 16'b0001110110010101;
            15'b001100011111101 : data = 16'b0001110110001000;
            15'b001100011111110 : data = 16'b0001110101111010;
            15'b001100011111111 : data = 16'b0001110101101101;
            15'b001100100000000 : data = 16'b0001110101100000;
            15'b001100100000001 : data = 16'b0001110101010011;
            15'b001100100000010 : data = 16'b0001110101000110;
            15'b001100100000011 : data = 16'b0001110100111001;
            15'b001100100000100 : data = 16'b0001110100101100;
            15'b001100100000101 : data = 16'b0001110100011111;
            15'b001100100000110 : data = 16'b0001110100010010;
            15'b001100100000111 : data = 16'b0001110100000100;
            15'b001100100001000 : data = 16'b0001110011110111;
            15'b001100100001001 : data = 16'b0001110011101010;
            15'b001100100001010 : data = 16'b0001110011011101;
            15'b001100100001011 : data = 16'b0001110011010000;
            15'b001100100001100 : data = 16'b0001110011000011;
            15'b001100100001101 : data = 16'b0001110010110110;
            15'b001100100001110 : data = 16'b0001110010101001;
            15'b001100100001111 : data = 16'b0001110010011100;
            15'b001100100010000 : data = 16'b0001110010001111;
            15'b001100100010001 : data = 16'b0001110010000010;
            15'b001100100010010 : data = 16'b0001110001110101;
            15'b001100100010011 : data = 16'b0001110001101001;
            15'b001100100010100 : data = 16'b0001110001011100;
            15'b001100100010101 : data = 16'b0001110001001111;
            15'b001100100010110 : data = 16'b0001110001000010;
            15'b001100100010111 : data = 16'b0001110000110101;
            15'b001100100011000 : data = 16'b0001110000101000;
            15'b001100100011001 : data = 16'b0001110000011011;
            15'b001100100011010 : data = 16'b0001110000001110;
            15'b001100100011011 : data = 16'b0001110000000001;
            15'b001100100011100 : data = 16'b0001101111110101;
            15'b001100100011101 : data = 16'b0001101111101000;
            15'b001100100011110 : data = 16'b0001101111011011;
            15'b001100100011111 : data = 16'b0001101111001110;
            15'b001100100100000 : data = 16'b0001101111000001;
            15'b001100100100001 : data = 16'b0001101110110100;
            15'b001100100100010 : data = 16'b0001101110101000;
            15'b001100100100011 : data = 16'b0001101110011011;
            15'b001100100100100 : data = 16'b0001101110001110;
            15'b001100100100101 : data = 16'b0001101110000001;
            15'b001100100100110 : data = 16'b0001101101110101;
            15'b001100100100111 : data = 16'b0001101101101000;
            15'b001100100101000 : data = 16'b0001101101011011;
            15'b001100100101001 : data = 16'b0001101101001110;
            15'b001100100101010 : data = 16'b0001101101000010;
            15'b001100100101011 : data = 16'b0001101100110101;
            15'b001100100101100 : data = 16'b0001101100101000;
            15'b001100100101101 : data = 16'b0001101100011100;
            15'b001100100101110 : data = 16'b0001101100001111;
            15'b001100100101111 : data = 16'b0001101100000010;
            15'b001100100110000 : data = 16'b0001101011110110;
            15'b001100100110001 : data = 16'b0001101011101001;
            15'b001100100110010 : data = 16'b0001101011011100;
            15'b001100100110011 : data = 16'b0001101011010000;
            15'b001100100110100 : data = 16'b0001101011000011;
            15'b001100100110101 : data = 16'b0001101010110111;
            15'b001100100110110 : data = 16'b0001101010101010;
            15'b001100100110111 : data = 16'b0001101010011110;
            15'b001100100111000 : data = 16'b0001101010010001;
            15'b001100100111001 : data = 16'b0001101010000100;
            15'b001100100111010 : data = 16'b0001101001111000;
            15'b001100100111011 : data = 16'b0001101001101011;
            15'b001100100111100 : data = 16'b0001101001011111;
            15'b001100100111101 : data = 16'b0001101001010010;
            15'b001100100111110 : data = 16'b0001101001000110;
            15'b001100100111111 : data = 16'b0001101000111001;
            15'b001100101000000 : data = 16'b0001101000101101;
            15'b001100101000001 : data = 16'b0001101000100000;
            15'b001100101000010 : data = 16'b0001101000010100;
            15'b001100101000011 : data = 16'b0001101000000111;
            15'b001100101000100 : data = 16'b0001100111111011;
            15'b001100101000101 : data = 16'b0001100111101111;
            15'b001100101000110 : data = 16'b0001100111100010;
            15'b001100101000111 : data = 16'b0001100111010110;
            15'b001100101001000 : data = 16'b0001100111001001;
            15'b001100101001001 : data = 16'b0001100110111101;
            15'b001100101001010 : data = 16'b0001100110110001;
            15'b001100101001011 : data = 16'b0001100110100100;
            15'b001100101001100 : data = 16'b0001100110011000;
            15'b001100101001101 : data = 16'b0001100110001100;
            15'b001100101001110 : data = 16'b0001100101111111;
            15'b001100101001111 : data = 16'b0001100101110011;
            15'b001100101010000 : data = 16'b0001100101100111;
            15'b001100101010001 : data = 16'b0001100101011010;
            15'b001100101010010 : data = 16'b0001100101001110;
            15'b001100101010011 : data = 16'b0001100101000010;
            15'b001100101010100 : data = 16'b0001100100110101;
            15'b001100101010101 : data = 16'b0001100100101001;
            15'b001100101010110 : data = 16'b0001100100011101;
            15'b001100101010111 : data = 16'b0001100100010001;
            15'b001100101011000 : data = 16'b0001100100000100;
            15'b001100101011001 : data = 16'b0001100011111000;
            15'b001100101011010 : data = 16'b0001100011101100;
            15'b001100101011011 : data = 16'b0001100011100000;
            15'b001100101011100 : data = 16'b0001100011010100;
            15'b001100101011101 : data = 16'b0001100011000111;
            15'b001100101011110 : data = 16'b0001100010111011;
            15'b001100101011111 : data = 16'b0001100010101111;
            15'b001100101100000 : data = 16'b0001100010100011;
            15'b001100101100001 : data = 16'b0001100010010111;
            15'b001100101100010 : data = 16'b0001100010001011;
            15'b001100101100011 : data = 16'b0001100001111111;
            15'b001100101100100 : data = 16'b0001100001110010;
            15'b001100101100101 : data = 16'b0001100001100110;
            15'b001100101100110 : data = 16'b0001100001011010;
            15'b001100101100111 : data = 16'b0001100001001110;
            15'b001100101101000 : data = 16'b0001100001000010;
            15'b001100101101001 : data = 16'b0001100000110110;
            15'b001100101101010 : data = 16'b0001100000101010;
            15'b001100101101011 : data = 16'b0001100000011110;
            15'b001100101101100 : data = 16'b0001100000010010;
            15'b001100101101101 : data = 16'b0001100000000110;
            15'b001100101101110 : data = 16'b0001011111111010;
            15'b001100101101111 : data = 16'b0001011111101110;
            15'b001100101110000 : data = 16'b0001011111100010;
            15'b001100101110001 : data = 16'b0001011111010110;
            15'b001100101110010 : data = 16'b0001011111001010;
            15'b001100101110011 : data = 16'b0001011110111110;
            15'b001100101110100 : data = 16'b0001011110110010;
            15'b001100101110101 : data = 16'b0001011110100110;
            15'b001100101110110 : data = 16'b0001011110011010;
            15'b001100101110111 : data = 16'b0001011110001110;
            15'b001100101111000 : data = 16'b0001011110000011;
            15'b001100101111001 : data = 16'b0001011101110111;
            15'b001100101111010 : data = 16'b0001011101101011;
            15'b001100101111011 : data = 16'b0001011101011111;
            15'b001100101111100 : data = 16'b0001011101010011;
            15'b001100101111101 : data = 16'b0001011101000111;
            15'b001100101111110 : data = 16'b0001011100111011;
            15'b001100101111111 : data = 16'b0001011100110000;
            15'b001100110000000 : data = 16'b0001011100100100;
            15'b001100110000001 : data = 16'b0001011100011000;
            15'b001100110000010 : data = 16'b0001011100001100;
            15'b001100110000011 : data = 16'b0001011100000000;
            15'b001100110000100 : data = 16'b0001011011110101;
            15'b001100110000101 : data = 16'b0001011011101001;
            15'b001100110000110 : data = 16'b0001011011011101;
            15'b001100110000111 : data = 16'b0001011011010001;
            15'b001100110001000 : data = 16'b0001011011000110;
            15'b001100110001001 : data = 16'b0001011010111010;
            15'b001100110001010 : data = 16'b0001011010101110;
            15'b001100110001011 : data = 16'b0001011010100010;
            15'b001100110001100 : data = 16'b0001011010010111;
            15'b001100110001101 : data = 16'b0001011010001011;
            15'b001100110001110 : data = 16'b0001011001111111;
            15'b001100110001111 : data = 16'b0001011001110100;
            15'b001100110010000 : data = 16'b0001011001101000;
            15'b001100110010001 : data = 16'b0001011001011101;
            15'b001100110010010 : data = 16'b0001011001010001;
            15'b001100110010011 : data = 16'b0001011001000101;
            15'b001100110010100 : data = 16'b0001011000111010;
            15'b001100110010101 : data = 16'b0001011000101110;
            15'b001100110010110 : data = 16'b0001011000100011;
            15'b001100110010111 : data = 16'b0001011000010111;
            15'b001100110011000 : data = 16'b0001011000001011;
            15'b001100110011001 : data = 16'b0001011000000000;
            15'b001100110011010 : data = 16'b0001010111110100;
            15'b001100110011011 : data = 16'b0001010111101001;
            15'b001100110011100 : data = 16'b0001010111011101;
            15'b001100110011101 : data = 16'b0001010111010010;
            15'b001100110011110 : data = 16'b0001010111000110;
            15'b001100110011111 : data = 16'b0001010110111011;
            15'b001100110100000 : data = 16'b0001010110101111;
            15'b001100110100001 : data = 16'b0001010110100100;
            15'b001100110100010 : data = 16'b0001010110011000;
            15'b001100110100011 : data = 16'b0001010110001101;
            15'b001100110100100 : data = 16'b0001010110000010;
            15'b001100110100101 : data = 16'b0001010101110110;
            15'b001100110100110 : data = 16'b0001010101101011;
            15'b001100110100111 : data = 16'b0001010101011111;
            15'b001100110101000 : data = 16'b0001010101010100;
            15'b001100110101001 : data = 16'b0001010101001001;
            15'b001100110101010 : data = 16'b0001010100111101;
            15'b001100110101011 : data = 16'b0001010100110010;
            15'b001100110101100 : data = 16'b0001010100100111;
            15'b001100110101101 : data = 16'b0001010100011011;
            15'b001100110101110 : data = 16'b0001010100010000;
            15'b001100110101111 : data = 16'b0001010100000101;
            15'b001100110110000 : data = 16'b0001010011111001;
            15'b001100110110001 : data = 16'b0001010011101110;
            15'b001100110110010 : data = 16'b0001010011100011;
            15'b001100110110011 : data = 16'b0001010011010111;
            15'b001100110110100 : data = 16'b0001010011001100;
            15'b001100110110101 : data = 16'b0001010011000001;
            15'b001100110110110 : data = 16'b0001010010110110;
            15'b001100110110111 : data = 16'b0001010010101011;
            15'b001100110111000 : data = 16'b0001010010011111;
            15'b001100110111001 : data = 16'b0001010010010100;
            15'b001100110111010 : data = 16'b0001010010001001;
            15'b001100110111011 : data = 16'b0001010001111110;
            15'b001100110111100 : data = 16'b0001010001110011;
            15'b001100110111101 : data = 16'b0001010001100111;
            15'b001100110111110 : data = 16'b0001010001011100;
            15'b001100110111111 : data = 16'b0001010001010001;
            15'b001100111000000 : data = 16'b0001010001000110;
            15'b001100111000001 : data = 16'b0001010000111011;
            15'b001100111000010 : data = 16'b0001010000110000;
            15'b001100111000011 : data = 16'b0001010000100101;
            15'b001100111000100 : data = 16'b0001010000011010;
            15'b001100111000101 : data = 16'b0001010000001111;
            15'b001100111000110 : data = 16'b0001010000000011;
            15'b001100111000111 : data = 16'b0001001111111000;
            15'b001100111001000 : data = 16'b0001001111101101;
            15'b001100111001001 : data = 16'b0001001111100010;
            15'b001100111001010 : data = 16'b0001001111010111;
            15'b001100111001011 : data = 16'b0001001111001100;
            15'b001100111001100 : data = 16'b0001001111000001;
            15'b001100111001101 : data = 16'b0001001110110110;
            15'b001100111001110 : data = 16'b0001001110101011;
            15'b001100111001111 : data = 16'b0001001110100000;
            15'b001100111010000 : data = 16'b0001001110010110;
            15'b001100111010001 : data = 16'b0001001110001011;
            15'b001100111010010 : data = 16'b0001001110000000;
            15'b001100111010011 : data = 16'b0001001101110101;
            15'b001100111010100 : data = 16'b0001001101101010;
            15'b001100111010101 : data = 16'b0001001101011111;
            15'b001100111010110 : data = 16'b0001001101010100;
            15'b001100111010111 : data = 16'b0001001101001001;
            15'b001100111011000 : data = 16'b0001001100111110;
            15'b001100111011001 : data = 16'b0001001100110011;
            15'b001100111011010 : data = 16'b0001001100101001;
            15'b001100111011011 : data = 16'b0001001100011110;
            15'b001100111011100 : data = 16'b0001001100010011;
            15'b001100111011101 : data = 16'b0001001100001000;
            15'b001100111011110 : data = 16'b0001001011111101;
            15'b001100111011111 : data = 16'b0001001011110011;
            15'b001100111100000 : data = 16'b0001001011101000;
            15'b001100111100001 : data = 16'b0001001011011101;
            15'b001100111100010 : data = 16'b0001001011010010;
            15'b001100111100011 : data = 16'b0001001011001000;
            15'b001100111100100 : data = 16'b0001001010111101;
            15'b001100111100101 : data = 16'b0001001010110010;
            15'b001100111100110 : data = 16'b0001001010100111;
            15'b001100111100111 : data = 16'b0001001010011101;
            15'b001100111101000 : data = 16'b0001001010010010;
            15'b001100111101001 : data = 16'b0001001010000111;
            15'b001100111101010 : data = 16'b0001001001111101;
            15'b001100111101011 : data = 16'b0001001001110010;
            15'b001100111101100 : data = 16'b0001001001100111;
            15'b001100111101101 : data = 16'b0001001001011101;
            15'b001100111101110 : data = 16'b0001001001010010;
            15'b001100111101111 : data = 16'b0001001001001000;
            15'b001100111110000 : data = 16'b0001001000111101;
            15'b001100111110001 : data = 16'b0001001000110010;
            15'b001100111110010 : data = 16'b0001001000101000;
            15'b001100111110011 : data = 16'b0001001000011101;
            15'b001100111110100 : data = 16'b0001001000010011;
            15'b001100111110101 : data = 16'b0001001000001000;
            15'b001100111110110 : data = 16'b0001000111111110;
            15'b001100111110111 : data = 16'b0001000111110011;
            15'b001100111111000 : data = 16'b0001000111101001;
            15'b001100111111001 : data = 16'b0001000111011110;
            15'b001100111111010 : data = 16'b0001000111010100;
            15'b001100111111011 : data = 16'b0001000111001001;
            15'b001100111111100 : data = 16'b0001000110111111;
            15'b001100111111101 : data = 16'b0001000110110100;
            15'b001100111111110 : data = 16'b0001000110101010;
            15'b001100111111111 : data = 16'b0001000110011111;
            15'b001101000000000 : data = 16'b0001000110010101;
            15'b001101000000001 : data = 16'b0001000110001010;
            15'b001101000000010 : data = 16'b0001000110000000;
            15'b001101000000011 : data = 16'b0001000101110110;
            15'b001101000000100 : data = 16'b0001000101101011;
            15'b001101000000101 : data = 16'b0001000101100001;
            15'b001101000000110 : data = 16'b0001000101010111;
            15'b001101000000111 : data = 16'b0001000101001100;
            15'b001101000001000 : data = 16'b0001000101000010;
            15'b001101000001001 : data = 16'b0001000100111000;
            15'b001101000001010 : data = 16'b0001000100101101;
            15'b001101000001011 : data = 16'b0001000100100011;
            15'b001101000001100 : data = 16'b0001000100011001;
            15'b001101000001101 : data = 16'b0001000100001110;
            15'b001101000001110 : data = 16'b0001000100000100;
            15'b001101000001111 : data = 16'b0001000011111010;
            15'b001101000010000 : data = 16'b0001000011110000;
            15'b001101000010001 : data = 16'b0001000011100101;
            15'b001101000010010 : data = 16'b0001000011011011;
            15'b001101000010011 : data = 16'b0001000011010001;
            15'b001101000010100 : data = 16'b0001000011000111;
            15'b001101000010101 : data = 16'b0001000010111101;
            15'b001101000010110 : data = 16'b0001000010110011;
            15'b001101000010111 : data = 16'b0001000010101000;
            15'b001101000011000 : data = 16'b0001000010011110;
            15'b001101000011001 : data = 16'b0001000010010100;
            15'b001101000011010 : data = 16'b0001000010001010;
            15'b001101000011011 : data = 16'b0001000010000000;
            15'b001101000011100 : data = 16'b0001000001110110;
            15'b001101000011101 : data = 16'b0001000001101100;
            15'b001101000011110 : data = 16'b0001000001100010;
            15'b001101000011111 : data = 16'b0001000001010111;
            15'b001101000100000 : data = 16'b0001000001001101;
            15'b001101000100001 : data = 16'b0001000001000011;
            15'b001101000100010 : data = 16'b0001000000111001;
            15'b001101000100011 : data = 16'b0001000000101111;
            15'b001101000100100 : data = 16'b0001000000100101;
            15'b001101000100101 : data = 16'b0001000000011011;
            15'b001101000100110 : data = 16'b0001000000010001;
            15'b001101000100111 : data = 16'b0001000000000111;
            15'b001101000101000 : data = 16'b0000111111111101;
            15'b001101000101001 : data = 16'b0000111111110011;
            15'b001101000101010 : data = 16'b0000111111101001;
            15'b001101000101011 : data = 16'b0000111111011111;
            15'b001101000101100 : data = 16'b0000111111010110;
            15'b001101000101101 : data = 16'b0000111111001100;
            15'b001101000101110 : data = 16'b0000111111000010;
            15'b001101000101111 : data = 16'b0000111110111000;
            15'b001101000110000 : data = 16'b0000111110101110;
            15'b001101000110001 : data = 16'b0000111110100100;
            15'b001101000110010 : data = 16'b0000111110011010;
            15'b001101000110011 : data = 16'b0000111110010000;
            15'b001101000110100 : data = 16'b0000111110000111;
            15'b001101000110101 : data = 16'b0000111101111101;
            15'b001101000110110 : data = 16'b0000111101110011;
            15'b001101000110111 : data = 16'b0000111101101001;
            15'b001101000111000 : data = 16'b0000111101011111;
            15'b001101000111001 : data = 16'b0000111101010110;
            15'b001101000111010 : data = 16'b0000111101001100;
            15'b001101000111011 : data = 16'b0000111101000010;
            15'b001101000111100 : data = 16'b0000111100111000;
            15'b001101000111101 : data = 16'b0000111100101111;
            15'b001101000111110 : data = 16'b0000111100100101;
            15'b001101000111111 : data = 16'b0000111100011011;
            15'b001101001000000 : data = 16'b0000111100010001;
            15'b001101001000001 : data = 16'b0000111100001000;
            15'b001101001000010 : data = 16'b0000111011111110;
            15'b001101001000011 : data = 16'b0000111011110100;
            15'b001101001000100 : data = 16'b0000111011101011;
            15'b001101001000101 : data = 16'b0000111011100001;
            15'b001101001000110 : data = 16'b0000111011011000;
            15'b001101001000111 : data = 16'b0000111011001110;
            15'b001101001001000 : data = 16'b0000111011000100;
            15'b001101001001001 : data = 16'b0000111010111011;
            15'b001101001001010 : data = 16'b0000111010110001;
            15'b001101001001011 : data = 16'b0000111010101000;
            15'b001101001001100 : data = 16'b0000111010011110;
            15'b001101001001101 : data = 16'b0000111010010100;
            15'b001101001001110 : data = 16'b0000111010001011;
            15'b001101001001111 : data = 16'b0000111010000001;
            15'b001101001010000 : data = 16'b0000111001111000;
            15'b001101001010001 : data = 16'b0000111001101110;
            15'b001101001010010 : data = 16'b0000111001100101;
            15'b001101001010011 : data = 16'b0000111001011011;
            15'b001101001010100 : data = 16'b0000111001010010;
            15'b001101001010101 : data = 16'b0000111001001000;
            15'b001101001010110 : data = 16'b0000111000111111;
            15'b001101001010111 : data = 16'b0000111000110110;
            15'b001101001011000 : data = 16'b0000111000101100;
            15'b001101001011001 : data = 16'b0000111000100011;
            15'b001101001011010 : data = 16'b0000111000011001;
            15'b001101001011011 : data = 16'b0000111000010000;
            15'b001101001011100 : data = 16'b0000111000000111;
            15'b001101001011101 : data = 16'b0000110111111101;
            15'b001101001011110 : data = 16'b0000110111110100;
            15'b001101001011111 : data = 16'b0000110111101011;
            15'b001101001100000 : data = 16'b0000110111100001;
            15'b001101001100001 : data = 16'b0000110111011000;
            15'b001101001100010 : data = 16'b0000110111001111;
            15'b001101001100011 : data = 16'b0000110111000101;
            15'b001101001100100 : data = 16'b0000110110111100;
            15'b001101001100101 : data = 16'b0000110110110011;
            15'b001101001100110 : data = 16'b0000110110101001;
            15'b001101001100111 : data = 16'b0000110110100000;
            15'b001101001101000 : data = 16'b0000110110010111;
            15'b001101001101001 : data = 16'b0000110110001110;
            15'b001101001101010 : data = 16'b0000110110000101;
            15'b001101001101011 : data = 16'b0000110101111011;
            15'b001101001101100 : data = 16'b0000110101110010;
            15'b001101001101101 : data = 16'b0000110101101001;
            15'b001101001101110 : data = 16'b0000110101100000;
            15'b001101001101111 : data = 16'b0000110101010111;
            15'b001101001110000 : data = 16'b0000110101001110;
            15'b001101001110001 : data = 16'b0000110101000100;
            15'b001101001110010 : data = 16'b0000110100111011;
            15'b001101001110011 : data = 16'b0000110100110010;
            15'b001101001110100 : data = 16'b0000110100101001;
            15'b001101001110101 : data = 16'b0000110100100000;
            15'b001101001110110 : data = 16'b0000110100010111;
            15'b001101001110111 : data = 16'b0000110100001110;
            15'b001101001111000 : data = 16'b0000110100000101;
            15'b001101001111001 : data = 16'b0000110011111100;
            15'b001101001111010 : data = 16'b0000110011110011;
            15'b001101001111011 : data = 16'b0000110011101010;
            15'b001101001111100 : data = 16'b0000110011100001;
            15'b001101001111101 : data = 16'b0000110011011000;
            15'b001101001111110 : data = 16'b0000110011001111;
            15'b001101001111111 : data = 16'b0000110011000110;
            15'b001101010000000 : data = 16'b0000110010111101;
            15'b001101010000001 : data = 16'b0000110010110100;
            15'b001101010000010 : data = 16'b0000110010101011;
            15'b001101010000011 : data = 16'b0000110010100010;
            15'b001101010000100 : data = 16'b0000110010011001;
            15'b001101010000101 : data = 16'b0000110010010000;
            15'b001101010000110 : data = 16'b0000110010000111;
            15'b001101010000111 : data = 16'b0000110001111110;
            15'b001101010001000 : data = 16'b0000110001110110;
            15'b001101010001001 : data = 16'b0000110001101101;
            15'b001101010001010 : data = 16'b0000110001100100;
            15'b001101010001011 : data = 16'b0000110001011011;
            15'b001101010001100 : data = 16'b0000110001010010;
            15'b001101010001101 : data = 16'b0000110001001001;
            15'b001101010001110 : data = 16'b0000110001000001;
            15'b001101010001111 : data = 16'b0000110000111000;
            15'b001101010010000 : data = 16'b0000110000101111;
            15'b001101010010001 : data = 16'b0000110000100110;
            15'b001101010010010 : data = 16'b0000110000011110;
            15'b001101010010011 : data = 16'b0000110000010101;
            15'b001101010010100 : data = 16'b0000110000001100;
            15'b001101010010101 : data = 16'b0000110000000011;
            15'b001101010010110 : data = 16'b0000101111111011;
            15'b001101010010111 : data = 16'b0000101111110010;
            15'b001101010011000 : data = 16'b0000101111101001;
            15'b001101010011001 : data = 16'b0000101111100001;
            15'b001101010011010 : data = 16'b0000101111011000;
            15'b001101010011011 : data = 16'b0000101111001111;
            15'b001101010011100 : data = 16'b0000101111000111;
            15'b001101010011101 : data = 16'b0000101110111110;
            15'b001101010011110 : data = 16'b0000101110110101;
            15'b001101010011111 : data = 16'b0000101110101101;
            15'b001101010100000 : data = 16'b0000101110100100;
            15'b001101010100001 : data = 16'b0000101110011100;
            15'b001101010100010 : data = 16'b0000101110010011;
            15'b001101010100011 : data = 16'b0000101110001011;
            15'b001101010100100 : data = 16'b0000101110000010;
            15'b001101010100101 : data = 16'b0000101101111010;
            15'b001101010100110 : data = 16'b0000101101110001;
            15'b001101010100111 : data = 16'b0000101101101001;
            15'b001101010101000 : data = 16'b0000101101100000;
            15'b001101010101001 : data = 16'b0000101101011000;
            15'b001101010101010 : data = 16'b0000101101001111;
            15'b001101010101011 : data = 16'b0000101101000111;
            15'b001101010101100 : data = 16'b0000101100111110;
            15'b001101010101101 : data = 16'b0000101100110110;
            15'b001101010101110 : data = 16'b0000101100101101;
            15'b001101010101111 : data = 16'b0000101100100101;
            15'b001101010110000 : data = 16'b0000101100011101;
            15'b001101010110001 : data = 16'b0000101100010100;
            15'b001101010110010 : data = 16'b0000101100001100;
            15'b001101010110011 : data = 16'b0000101100000011;
            15'b001101010110100 : data = 16'b0000101011111011;
            15'b001101010110101 : data = 16'b0000101011110011;
            15'b001101010110110 : data = 16'b0000101011101010;
            15'b001101010110111 : data = 16'b0000101011100010;
            15'b001101010111000 : data = 16'b0000101011011010;
            15'b001101010111001 : data = 16'b0000101011010010;
            15'b001101010111010 : data = 16'b0000101011001001;
            15'b001101010111011 : data = 16'b0000101011000001;
            15'b001101010111100 : data = 16'b0000101010111001;
            15'b001101010111101 : data = 16'b0000101010110000;
            15'b001101010111110 : data = 16'b0000101010101000;
            15'b001101010111111 : data = 16'b0000101010100000;
            15'b001101011000000 : data = 16'b0000101010011000;
            15'b001101011000001 : data = 16'b0000101010010000;
            15'b001101011000010 : data = 16'b0000101010000111;
            15'b001101011000011 : data = 16'b0000101001111111;
            15'b001101011000100 : data = 16'b0000101001110111;
            15'b001101011000101 : data = 16'b0000101001101111;
            15'b001101011000110 : data = 16'b0000101001100111;
            15'b001101011000111 : data = 16'b0000101001011111;
            15'b001101011001000 : data = 16'b0000101001010111;
            15'b001101011001001 : data = 16'b0000101001001110;
            15'b001101011001010 : data = 16'b0000101001000110;
            15'b001101011001011 : data = 16'b0000101000111110;
            15'b001101011001100 : data = 16'b0000101000110110;
            15'b001101011001101 : data = 16'b0000101000101110;
            15'b001101011001110 : data = 16'b0000101000100110;
            15'b001101011001111 : data = 16'b0000101000011110;
            15'b001101011010000 : data = 16'b0000101000010110;
            15'b001101011010001 : data = 16'b0000101000001110;
            15'b001101011010010 : data = 16'b0000101000000110;
            15'b001101011010011 : data = 16'b0000100111111110;
            15'b001101011010100 : data = 16'b0000100111110110;
            15'b001101011010101 : data = 16'b0000100111101110;
            15'b001101011010110 : data = 16'b0000100111100110;
            15'b001101011010111 : data = 16'b0000100111011110;
            15'b001101011011000 : data = 16'b0000100111010110;
            15'b001101011011001 : data = 16'b0000100111001111;
            15'b001101011011010 : data = 16'b0000100111000111;
            15'b001101011011011 : data = 16'b0000100110111111;
            15'b001101011011100 : data = 16'b0000100110110111;
            15'b001101011011101 : data = 16'b0000100110101111;
            15'b001101011011110 : data = 16'b0000100110100111;
            15'b001101011011111 : data = 16'b0000100110011111;
            15'b001101011100000 : data = 16'b0000100110010111;
            15'b001101011100001 : data = 16'b0000100110010000;
            15'b001101011100010 : data = 16'b0000100110001000;
            15'b001101011100011 : data = 16'b0000100110000000;
            15'b001101011100100 : data = 16'b0000100101111000;
            15'b001101011100101 : data = 16'b0000100101110001;
            15'b001101011100110 : data = 16'b0000100101101001;
            15'b001101011100111 : data = 16'b0000100101100001;
            15'b001101011101000 : data = 16'b0000100101011001;
            15'b001101011101001 : data = 16'b0000100101010010;
            15'b001101011101010 : data = 16'b0000100101001010;
            15'b001101011101011 : data = 16'b0000100101000010;
            15'b001101011101100 : data = 16'b0000100100111011;
            15'b001101011101101 : data = 16'b0000100100110011;
            15'b001101011101110 : data = 16'b0000100100101011;
            15'b001101011101111 : data = 16'b0000100100100100;
            15'b001101011110000 : data = 16'b0000100100011100;
            15'b001101011110001 : data = 16'b0000100100010100;
            15'b001101011110010 : data = 16'b0000100100001101;
            15'b001101011110011 : data = 16'b0000100100000101;
            15'b001101011110100 : data = 16'b0000100011111110;
            15'b001101011110101 : data = 16'b0000100011110110;
            15'b001101011110110 : data = 16'b0000100011101110;
            15'b001101011110111 : data = 16'b0000100011100111;
            15'b001101011111000 : data = 16'b0000100011011111;
            15'b001101011111001 : data = 16'b0000100011011000;
            15'b001101011111010 : data = 16'b0000100011010000;
            15'b001101011111011 : data = 16'b0000100011001001;
            15'b001101011111100 : data = 16'b0000100011000001;
            15'b001101011111101 : data = 16'b0000100010111010;
            15'b001101011111110 : data = 16'b0000100010110010;
            15'b001101011111111 : data = 16'b0000100010101011;
            15'b001101100000000 : data = 16'b0000100010100011;
            15'b001101100000001 : data = 16'b0000100010011100;
            15'b001101100000010 : data = 16'b0000100010010101;
            15'b001101100000011 : data = 16'b0000100010001101;
            15'b001101100000100 : data = 16'b0000100010000110;
            15'b001101100000101 : data = 16'b0000100001111110;
            15'b001101100000110 : data = 16'b0000100001110111;
            15'b001101100000111 : data = 16'b0000100001110000;
            15'b001101100001000 : data = 16'b0000100001101000;
            15'b001101100001001 : data = 16'b0000100001100001;
            15'b001101100001010 : data = 16'b0000100001011010;
            15'b001101100001011 : data = 16'b0000100001010010;
            15'b001101100001100 : data = 16'b0000100001001011;
            15'b001101100001101 : data = 16'b0000100001000100;
            15'b001101100001110 : data = 16'b0000100000111101;
            15'b001101100001111 : data = 16'b0000100000110101;
            15'b001101100010000 : data = 16'b0000100000101110;
            15'b001101100010001 : data = 16'b0000100000100111;
            15'b001101100010010 : data = 16'b0000100000100000;
            15'b001101100010011 : data = 16'b0000100000011000;
            15'b001101100010100 : data = 16'b0000100000010001;
            15'b001101100010101 : data = 16'b0000100000001010;
            15'b001101100010110 : data = 16'b0000100000000011;
            15'b001101100010111 : data = 16'b0000011111111100;
            15'b001101100011000 : data = 16'b0000011111110100;
            15'b001101100011001 : data = 16'b0000011111101101;
            15'b001101100011010 : data = 16'b0000011111100110;
            15'b001101100011011 : data = 16'b0000011111011111;
            15'b001101100011100 : data = 16'b0000011111011000;
            15'b001101100011101 : data = 16'b0000011111010001;
            15'b001101100011110 : data = 16'b0000011111001010;
            15'b001101100011111 : data = 16'b0000011111000011;
            15'b001101100100000 : data = 16'b0000011110111100;
            15'b001101100100001 : data = 16'b0000011110110101;
            15'b001101100100010 : data = 16'b0000011110101110;
            15'b001101100100011 : data = 16'b0000011110100111;
            15'b001101100100100 : data = 16'b0000011110100000;
            15'b001101100100101 : data = 16'b0000011110011001;
            15'b001101100100110 : data = 16'b0000011110010010;
            15'b001101100100111 : data = 16'b0000011110001011;
            15'b001101100101000 : data = 16'b0000011110000100;
            15'b001101100101001 : data = 16'b0000011101111101;
            15'b001101100101010 : data = 16'b0000011101110110;
            15'b001101100101011 : data = 16'b0000011101101111;
            15'b001101100101100 : data = 16'b0000011101101000;
            15'b001101100101101 : data = 16'b0000011101100001;
            15'b001101100101110 : data = 16'b0000011101011010;
            15'b001101100101111 : data = 16'b0000011101010011;
            15'b001101100110000 : data = 16'b0000011101001101;
            15'b001101100110001 : data = 16'b0000011101000110;
            15'b001101100110010 : data = 16'b0000011100111111;
            15'b001101100110011 : data = 16'b0000011100111000;
            15'b001101100110100 : data = 16'b0000011100110001;
            15'b001101100110101 : data = 16'b0000011100101010;
            15'b001101100110110 : data = 16'b0000011100100100;
            15'b001101100110111 : data = 16'b0000011100011101;
            15'b001101100111000 : data = 16'b0000011100010110;
            15'b001101100111001 : data = 16'b0000011100001111;
            15'b001101100111010 : data = 16'b0000011100001001;
            15'b001101100111011 : data = 16'b0000011100000010;
            15'b001101100111100 : data = 16'b0000011011111011;
            15'b001101100111101 : data = 16'b0000011011110100;
            15'b001101100111110 : data = 16'b0000011011101110;
            15'b001101100111111 : data = 16'b0000011011100111;
            15'b001101101000000 : data = 16'b0000011011100000;
            15'b001101101000001 : data = 16'b0000011011011010;
            15'b001101101000010 : data = 16'b0000011011010011;
            15'b001101101000011 : data = 16'b0000011011001101;
            15'b001101101000100 : data = 16'b0000011011000110;
            15'b001101101000101 : data = 16'b0000011010111111;
            15'b001101101000110 : data = 16'b0000011010111001;
            15'b001101101000111 : data = 16'b0000011010110010;
            15'b001101101001000 : data = 16'b0000011010101100;
            15'b001101101001001 : data = 16'b0000011010100101;
            15'b001101101001010 : data = 16'b0000011010011111;
            15'b001101101001011 : data = 16'b0000011010011000;
            15'b001101101001100 : data = 16'b0000011010010001;
            15'b001101101001101 : data = 16'b0000011010001011;
            15'b001101101001110 : data = 16'b0000011010000100;
            15'b001101101001111 : data = 16'b0000011001111110;
            15'b001101101010000 : data = 16'b0000011001111000;
            15'b001101101010001 : data = 16'b0000011001110001;
            15'b001101101010010 : data = 16'b0000011001101011;
            15'b001101101010011 : data = 16'b0000011001100100;
            15'b001101101010100 : data = 16'b0000011001011110;
            15'b001101101010101 : data = 16'b0000011001010111;
            15'b001101101010110 : data = 16'b0000011001010001;
            15'b001101101010111 : data = 16'b0000011001001011;
            15'b001101101011000 : data = 16'b0000011001000100;
            15'b001101101011001 : data = 16'b0000011000111110;
            15'b001101101011010 : data = 16'b0000011000111000;
            15'b001101101011011 : data = 16'b0000011000110001;
            15'b001101101011100 : data = 16'b0000011000101011;
            15'b001101101011101 : data = 16'b0000011000100101;
            15'b001101101011110 : data = 16'b0000011000011110;
            15'b001101101011111 : data = 16'b0000011000011000;
            15'b001101101100000 : data = 16'b0000011000010010;
            15'b001101101100001 : data = 16'b0000011000001011;
            15'b001101101100010 : data = 16'b0000011000000101;
            15'b001101101100011 : data = 16'b0000010111111111;
            15'b001101101100100 : data = 16'b0000010111111001;
            15'b001101101100101 : data = 16'b0000010111110011;
            15'b001101101100110 : data = 16'b0000010111101100;
            15'b001101101100111 : data = 16'b0000010111100110;
            15'b001101101101000 : data = 16'b0000010111100000;
            15'b001101101101001 : data = 16'b0000010111011010;
            15'b001101101101010 : data = 16'b0000010111010100;
            15'b001101101101011 : data = 16'b0000010111001110;
            15'b001101101101100 : data = 16'b0000010111000111;
            15'b001101101101101 : data = 16'b0000010111000001;
            15'b001101101101110 : data = 16'b0000010110111011;
            15'b001101101101111 : data = 16'b0000010110110101;
            15'b001101101110000 : data = 16'b0000010110101111;
            15'b001101101110001 : data = 16'b0000010110101001;
            15'b001101101110010 : data = 16'b0000010110100011;
            15'b001101101110011 : data = 16'b0000010110011101;
            15'b001101101110100 : data = 16'b0000010110010111;
            15'b001101101110101 : data = 16'b0000010110010001;
            15'b001101101110110 : data = 16'b0000010110001011;
            15'b001101101110111 : data = 16'b0000010110000101;
            15'b001101101111000 : data = 16'b0000010101111111;
            15'b001101101111001 : data = 16'b0000010101111001;
            15'b001101101111010 : data = 16'b0000010101110011;
            15'b001101101111011 : data = 16'b0000010101101101;
            15'b001101101111100 : data = 16'b0000010101100111;
            15'b001101101111101 : data = 16'b0000010101100001;
            15'b001101101111110 : data = 16'b0000010101011011;
            15'b001101101111111 : data = 16'b0000010101010101;
            15'b001101110000000 : data = 16'b0000010101010000;
            15'b001101110000001 : data = 16'b0000010101001010;
            15'b001101110000010 : data = 16'b0000010101000100;
            15'b001101110000011 : data = 16'b0000010100111110;
            15'b001101110000100 : data = 16'b0000010100111000;
            15'b001101110000101 : data = 16'b0000010100110010;
            15'b001101110000110 : data = 16'b0000010100101101;
            15'b001101110000111 : data = 16'b0000010100100111;
            15'b001101110001000 : data = 16'b0000010100100001;
            15'b001101110001001 : data = 16'b0000010100011011;
            15'b001101110001010 : data = 16'b0000010100010110;
            15'b001101110001011 : data = 16'b0000010100010000;
            15'b001101110001100 : data = 16'b0000010100001010;
            15'b001101110001101 : data = 16'b0000010100000100;
            15'b001101110001110 : data = 16'b0000010011111111;
            15'b001101110001111 : data = 16'b0000010011111001;
            15'b001101110010000 : data = 16'b0000010011110011;
            15'b001101110010001 : data = 16'b0000010011101110;
            15'b001101110010010 : data = 16'b0000010011101000;
            15'b001101110010011 : data = 16'b0000010011100010;
            15'b001101110010100 : data = 16'b0000010011011101;
            15'b001101110010101 : data = 16'b0000010011010111;
            15'b001101110010110 : data = 16'b0000010011010010;
            15'b001101110010111 : data = 16'b0000010011001100;
            15'b001101110011000 : data = 16'b0000010011000110;
            15'b001101110011001 : data = 16'b0000010011000001;
            15'b001101110011010 : data = 16'b0000010010111011;
            15'b001101110011011 : data = 16'b0000010010110110;
            15'b001101110011100 : data = 16'b0000010010110000;
            15'b001101110011101 : data = 16'b0000010010101011;
            15'b001101110011110 : data = 16'b0000010010100101;
            15'b001101110011111 : data = 16'b0000010010100000;
            15'b001101110100000 : data = 16'b0000010010011010;
            15'b001101110100001 : data = 16'b0000010010010101;
            15'b001101110100010 : data = 16'b0000010010001111;
            15'b001101110100011 : data = 16'b0000010010001010;
            15'b001101110100100 : data = 16'b0000010010000100;
            15'b001101110100101 : data = 16'b0000010001111111;
            15'b001101110100110 : data = 16'b0000010001111010;
            15'b001101110100111 : data = 16'b0000010001110100;
            15'b001101110101000 : data = 16'b0000010001101111;
            15'b001101110101001 : data = 16'b0000010001101001;
            15'b001101110101010 : data = 16'b0000010001100100;
            15'b001101110101011 : data = 16'b0000010001011111;
            15'b001101110101100 : data = 16'b0000010001011001;
            15'b001101110101101 : data = 16'b0000010001010100;
            15'b001101110101110 : data = 16'b0000010001001111;
            15'b001101110101111 : data = 16'b0000010001001010;
            15'b001101110110000 : data = 16'b0000010001000100;
            15'b001101110110001 : data = 16'b0000010000111111;
            15'b001101110110010 : data = 16'b0000010000111010;
            15'b001101110110011 : data = 16'b0000010000110101;
            15'b001101110110100 : data = 16'b0000010000101111;
            15'b001101110110101 : data = 16'b0000010000101010;
            15'b001101110110110 : data = 16'b0000010000100101;
            15'b001101110110111 : data = 16'b0000010000100000;
            15'b001101110111000 : data = 16'b0000010000011011;
            15'b001101110111001 : data = 16'b0000010000010101;
            15'b001101110111010 : data = 16'b0000010000010000;
            15'b001101110111011 : data = 16'b0000010000001011;
            15'b001101110111100 : data = 16'b0000010000000110;
            15'b001101110111101 : data = 16'b0000010000000001;
            15'b001101110111110 : data = 16'b0000001111111100;
            15'b001101110111111 : data = 16'b0000001111110111;
            15'b001101111000000 : data = 16'b0000001111110010;
            15'b001101111000001 : data = 16'b0000001111101100;
            15'b001101111000010 : data = 16'b0000001111100111;
            15'b001101111000011 : data = 16'b0000001111100010;
            15'b001101111000100 : data = 16'b0000001111011101;
            15'b001101111000101 : data = 16'b0000001111011000;
            15'b001101111000110 : data = 16'b0000001111010011;
            15'b001101111000111 : data = 16'b0000001111001110;
            15'b001101111001000 : data = 16'b0000001111001001;
            15'b001101111001001 : data = 16'b0000001111000100;
            15'b001101111001010 : data = 16'b0000001110111111;
            15'b001101111001011 : data = 16'b0000001110111011;
            15'b001101111001100 : data = 16'b0000001110110110;
            15'b001101111001101 : data = 16'b0000001110110001;
            15'b001101111001110 : data = 16'b0000001110101100;
            15'b001101111001111 : data = 16'b0000001110100111;
            15'b001101111010000 : data = 16'b0000001110100010;
            15'b001101111010001 : data = 16'b0000001110011101;
            15'b001101111010010 : data = 16'b0000001110011000;
            15'b001101111010011 : data = 16'b0000001110010011;
            15'b001101111010100 : data = 16'b0000001110001111;
            15'b001101111010101 : data = 16'b0000001110001010;
            15'b001101111010110 : data = 16'b0000001110000101;
            15'b001101111010111 : data = 16'b0000001110000000;
            15'b001101111011000 : data = 16'b0000001101111011;
            15'b001101111011001 : data = 16'b0000001101110111;
            15'b001101111011010 : data = 16'b0000001101110010;
            15'b001101111011011 : data = 16'b0000001101101101;
            15'b001101111011100 : data = 16'b0000001101101001;
            15'b001101111011101 : data = 16'b0000001101100100;
            15'b001101111011110 : data = 16'b0000001101011111;
            15'b001101111011111 : data = 16'b0000001101011010;
            15'b001101111100000 : data = 16'b0000001101010110;
            15'b001101111100001 : data = 16'b0000001101010001;
            15'b001101111100010 : data = 16'b0000001101001100;
            15'b001101111100011 : data = 16'b0000001101001000;
            15'b001101111100100 : data = 16'b0000001101000011;
            15'b001101111100101 : data = 16'b0000001100111111;
            15'b001101111100110 : data = 16'b0000001100111010;
            15'b001101111100111 : data = 16'b0000001100110101;
            15'b001101111101000 : data = 16'b0000001100110001;
            15'b001101111101001 : data = 16'b0000001100101100;
            15'b001101111101010 : data = 16'b0000001100101000;
            15'b001101111101011 : data = 16'b0000001100100011;
            15'b001101111101100 : data = 16'b0000001100011111;
            15'b001101111101101 : data = 16'b0000001100011010;
            15'b001101111101110 : data = 16'b0000001100010110;
            15'b001101111101111 : data = 16'b0000001100010001;
            15'b001101111110000 : data = 16'b0000001100001101;
            15'b001101111110001 : data = 16'b0000001100001000;
            15'b001101111110010 : data = 16'b0000001100000100;
            15'b001101111110011 : data = 16'b0000001011111111;
            15'b001101111110100 : data = 16'b0000001011111011;
            15'b001101111110101 : data = 16'b0000001011110111;
            15'b001101111110110 : data = 16'b0000001011110010;
            15'b001101111110111 : data = 16'b0000001011101110;
            15'b001101111111000 : data = 16'b0000001011101001;
            15'b001101111111001 : data = 16'b0000001011100101;
            15'b001101111111010 : data = 16'b0000001011100001;
            15'b001101111111011 : data = 16'b0000001011011100;
            15'b001101111111100 : data = 16'b0000001011011000;
            15'b001101111111101 : data = 16'b0000001011010100;
            15'b001101111111110 : data = 16'b0000001011001111;
            15'b001101111111111 : data = 16'b0000001011001011;
            15'b001110000000000 : data = 16'b0000001011000111;
            15'b001110000000001 : data = 16'b0000001011000011;
            15'b001110000000010 : data = 16'b0000001010111110;
            15'b001110000000011 : data = 16'b0000001010111010;
            15'b001110000000100 : data = 16'b0000001010110110;
            15'b001110000000101 : data = 16'b0000001010110010;
            15'b001110000000110 : data = 16'b0000001010101101;
            15'b001110000000111 : data = 16'b0000001010101001;
            15'b001110000001000 : data = 16'b0000001010100101;
            15'b001110000001001 : data = 16'b0000001010100001;
            15'b001110000001010 : data = 16'b0000001010011101;
            15'b001110000001011 : data = 16'b0000001010011001;
            15'b001110000001100 : data = 16'b0000001010010101;
            15'b001110000001101 : data = 16'b0000001010010000;
            15'b001110000001110 : data = 16'b0000001010001100;
            15'b001110000001111 : data = 16'b0000001010001000;
            15'b001110000010000 : data = 16'b0000001010000100;
            15'b001110000010001 : data = 16'b0000001010000000;
            15'b001110000010010 : data = 16'b0000001001111100;
            15'b001110000010011 : data = 16'b0000001001111000;
            15'b001110000010100 : data = 16'b0000001001110100;
            15'b001110000010101 : data = 16'b0000001001110000;
            15'b001110000010110 : data = 16'b0000001001101100;
            15'b001110000010111 : data = 16'b0000001001101000;
            15'b001110000011000 : data = 16'b0000001001100100;
            15'b001110000011001 : data = 16'b0000001001100000;
            15'b001110000011010 : data = 16'b0000001001011100;
            15'b001110000011011 : data = 16'b0000001001011000;
            15'b001110000011100 : data = 16'b0000001001010100;
            15'b001110000011101 : data = 16'b0000001001010001;
            15'b001110000011110 : data = 16'b0000001001001101;
            15'b001110000011111 : data = 16'b0000001001001001;
            15'b001110000100000 : data = 16'b0000001001000101;
            15'b001110000100001 : data = 16'b0000001001000001;
            15'b001110000100010 : data = 16'b0000001000111101;
            15'b001110000100011 : data = 16'b0000001000111001;
            15'b001110000100100 : data = 16'b0000001000110110;
            15'b001110000100101 : data = 16'b0000001000110010;
            15'b001110000100110 : data = 16'b0000001000101110;
            15'b001110000100111 : data = 16'b0000001000101010;
            15'b001110000101000 : data = 16'b0000001000100110;
            15'b001110000101001 : data = 16'b0000001000100011;
            15'b001110000101010 : data = 16'b0000001000011111;
            15'b001110000101011 : data = 16'b0000001000011011;
            15'b001110000101100 : data = 16'b0000001000011000;
            15'b001110000101101 : data = 16'b0000001000010100;
            15'b001110000101110 : data = 16'b0000001000010000;
            15'b001110000101111 : data = 16'b0000001000001100;
            15'b001110000110000 : data = 16'b0000001000001001;
            15'b001110000110001 : data = 16'b0000001000000101;
            15'b001110000110010 : data = 16'b0000001000000010;
            15'b001110000110011 : data = 16'b0000000111111110;
            15'b001110000110100 : data = 16'b0000000111111010;
            15'b001110000110101 : data = 16'b0000000111110111;
            15'b001110000110110 : data = 16'b0000000111110011;
            15'b001110000110111 : data = 16'b0000000111110000;
            15'b001110000111000 : data = 16'b0000000111101100;
            15'b001110000111001 : data = 16'b0000000111101000;
            15'b001110000111010 : data = 16'b0000000111100101;
            15'b001110000111011 : data = 16'b0000000111100001;
            15'b001110000111100 : data = 16'b0000000111011110;
            15'b001110000111101 : data = 16'b0000000111011010;
            15'b001110000111110 : data = 16'b0000000111010111;
            15'b001110000111111 : data = 16'b0000000111010011;
            15'b001110001000000 : data = 16'b0000000111010000;
            15'b001110001000001 : data = 16'b0000000111001101;
            15'b001110001000010 : data = 16'b0000000111001001;
            15'b001110001000011 : data = 16'b0000000111000110;
            15'b001110001000100 : data = 16'b0000000111000010;
            15'b001110001000101 : data = 16'b0000000110111111;
            15'b001110001000110 : data = 16'b0000000110111011;
            15'b001110001000111 : data = 16'b0000000110111000;
            15'b001110001001000 : data = 16'b0000000110110101;
            15'b001110001001001 : data = 16'b0000000110110001;
            15'b001110001001010 : data = 16'b0000000110101110;
            15'b001110001001011 : data = 16'b0000000110101011;
            15'b001110001001100 : data = 16'b0000000110100111;
            15'b001110001001101 : data = 16'b0000000110100100;
            15'b001110001001110 : data = 16'b0000000110100001;
            15'b001110001001111 : data = 16'b0000000110011110;
            15'b001110001010000 : data = 16'b0000000110011010;
            15'b001110001010001 : data = 16'b0000000110010111;
            15'b001110001010010 : data = 16'b0000000110010100;
            15'b001110001010011 : data = 16'b0000000110010001;
            15'b001110001010100 : data = 16'b0000000110001110;
            15'b001110001010101 : data = 16'b0000000110001010;
            15'b001110001010110 : data = 16'b0000000110000111;
            15'b001110001010111 : data = 16'b0000000110000100;
            15'b001110001011000 : data = 16'b0000000110000001;
            15'b001110001011001 : data = 16'b0000000101111110;
            15'b001110001011010 : data = 16'b0000000101111011;
            15'b001110001011011 : data = 16'b0000000101110111;
            15'b001110001011100 : data = 16'b0000000101110100;
            15'b001110001011101 : data = 16'b0000000101110001;
            15'b001110001011110 : data = 16'b0000000101101110;
            15'b001110001011111 : data = 16'b0000000101101011;
            15'b001110001100000 : data = 16'b0000000101101000;
            15'b001110001100001 : data = 16'b0000000101100101;
            15'b001110001100010 : data = 16'b0000000101100010;
            15'b001110001100011 : data = 16'b0000000101011111;
            15'b001110001100100 : data = 16'b0000000101011100;
            15'b001110001100101 : data = 16'b0000000101011001;
            15'b001110001100110 : data = 16'b0000000101010110;
            15'b001110001100111 : data = 16'b0000000101010011;
            15'b001110001101000 : data = 16'b0000000101010000;
            15'b001110001101001 : data = 16'b0000000101001101;
            15'b001110001101010 : data = 16'b0000000101001010;
            15'b001110001101011 : data = 16'b0000000101000111;
            15'b001110001101100 : data = 16'b0000000101000101;
            15'b001110001101101 : data = 16'b0000000101000010;
            15'b001110001101110 : data = 16'b0000000100111111;
            15'b001110001101111 : data = 16'b0000000100111100;
            15'b001110001110000 : data = 16'b0000000100111001;
            15'b001110001110001 : data = 16'b0000000100110110;
            15'b001110001110010 : data = 16'b0000000100110011;
            15'b001110001110011 : data = 16'b0000000100110001;
            15'b001110001110100 : data = 16'b0000000100101110;
            15'b001110001110101 : data = 16'b0000000100101011;
            15'b001110001110110 : data = 16'b0000000100101000;
            15'b001110001110111 : data = 16'b0000000100100110;
            15'b001110001111000 : data = 16'b0000000100100011;
            15'b001110001111001 : data = 16'b0000000100100000;
            15'b001110001111010 : data = 16'b0000000100011101;
            15'b001110001111011 : data = 16'b0000000100011011;
            15'b001110001111100 : data = 16'b0000000100011000;
            15'b001110001111101 : data = 16'b0000000100010101;
            15'b001110001111110 : data = 16'b0000000100010011;
            15'b001110001111111 : data = 16'b0000000100010000;
            15'b001110010000000 : data = 16'b0000000100001101;
            15'b001110010000001 : data = 16'b0000000100001011;
            15'b001110010000010 : data = 16'b0000000100001000;
            15'b001110010000011 : data = 16'b0000000100000101;
            15'b001110010000100 : data = 16'b0000000100000011;
            15'b001110010000101 : data = 16'b0000000100000000;
            15'b001110010000110 : data = 16'b0000000011111110;
            15'b001110010000111 : data = 16'b0000000011111011;
            15'b001110010001000 : data = 16'b0000000011111001;
            15'b001110010001001 : data = 16'b0000000011110110;
            15'b001110010001010 : data = 16'b0000000011110100;
            15'b001110010001011 : data = 16'b0000000011110001;
            15'b001110010001100 : data = 16'b0000000011101111;
            15'b001110010001101 : data = 16'b0000000011101100;
            15'b001110010001110 : data = 16'b0000000011101010;
            15'b001110010001111 : data = 16'b0000000011100111;
            15'b001110010010000 : data = 16'b0000000011100101;
            15'b001110010010001 : data = 16'b0000000011100010;
            15'b001110010010010 : data = 16'b0000000011100000;
            15'b001110010010011 : data = 16'b0000000011011110;
            15'b001110010010100 : data = 16'b0000000011011011;
            15'b001110010010101 : data = 16'b0000000011011001;
            15'b001110010010110 : data = 16'b0000000011010111;
            15'b001110010010111 : data = 16'b0000000011010100;
            15'b001110010011000 : data = 16'b0000000011010010;
            15'b001110010011001 : data = 16'b0000000011010000;
            15'b001110010011010 : data = 16'b0000000011001101;
            15'b001110010011011 : data = 16'b0000000011001011;
            15'b001110010011100 : data = 16'b0000000011001001;
            15'b001110010011101 : data = 16'b0000000011000110;
            15'b001110010011110 : data = 16'b0000000011000100;
            15'b001110010011111 : data = 16'b0000000011000010;
            15'b001110010100000 : data = 16'b0000000011000000;
            15'b001110010100001 : data = 16'b0000000010111101;
            15'b001110010100010 : data = 16'b0000000010111011;
            15'b001110010100011 : data = 16'b0000000010111001;
            15'b001110010100100 : data = 16'b0000000010110111;
            15'b001110010100101 : data = 16'b0000000010110101;
            15'b001110010100110 : data = 16'b0000000010110011;
            15'b001110010100111 : data = 16'b0000000010110000;
            15'b001110010101000 : data = 16'b0000000010101110;
            15'b001110010101001 : data = 16'b0000000010101100;
            15'b001110010101010 : data = 16'b0000000010101010;
            15'b001110010101011 : data = 16'b0000000010101000;
            15'b001110010101100 : data = 16'b0000000010100110;
            15'b001110010101101 : data = 16'b0000000010100100;
            15'b001110010101110 : data = 16'b0000000010100010;
            15'b001110010101111 : data = 16'b0000000010100000;
            15'b001110010110000 : data = 16'b0000000010011110;
            15'b001110010110001 : data = 16'b0000000010011100;
            15'b001110010110010 : data = 16'b0000000010011010;
            15'b001110010110011 : data = 16'b0000000010011000;
            15'b001110010110100 : data = 16'b0000000010010110;
            15'b001110010110101 : data = 16'b0000000010010100;
            15'b001110010110110 : data = 16'b0000000010010010;
            15'b001110010110111 : data = 16'b0000000010010000;
            15'b001110010111000 : data = 16'b0000000010001110;
            15'b001110010111001 : data = 16'b0000000010001100;
            15'b001110010111010 : data = 16'b0000000010001010;
            15'b001110010111011 : data = 16'b0000000010001000;
            15'b001110010111100 : data = 16'b0000000010000111;
            15'b001110010111101 : data = 16'b0000000010000101;
            15'b001110010111110 : data = 16'b0000000010000011;
            15'b001110010111111 : data = 16'b0000000010000001;
            15'b001110011000000 : data = 16'b0000000001111111;
            15'b001110011000001 : data = 16'b0000000001111101;
            15'b001110011000010 : data = 16'b0000000001111100;
            15'b001110011000011 : data = 16'b0000000001111010;
            15'b001110011000100 : data = 16'b0000000001111000;
            15'b001110011000101 : data = 16'b0000000001110110;
            15'b001110011000110 : data = 16'b0000000001110101;
            15'b001110011000111 : data = 16'b0000000001110011;
            15'b001110011001000 : data = 16'b0000000001110001;
            15'b001110011001001 : data = 16'b0000000001101111;
            15'b001110011001010 : data = 16'b0000000001101110;
            15'b001110011001011 : data = 16'b0000000001101100;
            15'b001110011001100 : data = 16'b0000000001101010;
            15'b001110011001101 : data = 16'b0000000001101001;
            15'b001110011001110 : data = 16'b0000000001100111;
            15'b001110011001111 : data = 16'b0000000001100110;
            15'b001110011010000 : data = 16'b0000000001100100;
            15'b001110011010001 : data = 16'b0000000001100010;
            15'b001110011010010 : data = 16'b0000000001100001;
            15'b001110011010011 : data = 16'b0000000001011111;
            15'b001110011010100 : data = 16'b0000000001011110;
            15'b001110011010101 : data = 16'b0000000001011100;
            15'b001110011010110 : data = 16'b0000000001011011;
            15'b001110011010111 : data = 16'b0000000001011001;
            15'b001110011011000 : data = 16'b0000000001010111;
            15'b001110011011001 : data = 16'b0000000001010110;
            15'b001110011011010 : data = 16'b0000000001010101;
            15'b001110011011011 : data = 16'b0000000001010011;
            15'b001110011011100 : data = 16'b0000000001010010;
            15'b001110011011101 : data = 16'b0000000001010000;
            15'b001110011011110 : data = 16'b0000000001001111;
            15'b001110011011111 : data = 16'b0000000001001101;
            15'b001110011100000 : data = 16'b0000000001001100;
            15'b001110011100001 : data = 16'b0000000001001011;
            15'b001110011100010 : data = 16'b0000000001001001;
            15'b001110011100011 : data = 16'b0000000001001000;
            15'b001110011100100 : data = 16'b0000000001000110;
            15'b001110011100101 : data = 16'b0000000001000101;
            15'b001110011100110 : data = 16'b0000000001000100;
            15'b001110011100111 : data = 16'b0000000001000010;
            15'b001110011101000 : data = 16'b0000000001000001;
            15'b001110011101001 : data = 16'b0000000001000000;
            15'b001110011101010 : data = 16'b0000000000111111;
            15'b001110011101011 : data = 16'b0000000000111101;
            15'b001110011101100 : data = 16'b0000000000111100;
            15'b001110011101101 : data = 16'b0000000000111011;
            15'b001110011101110 : data = 16'b0000000000111010;
            15'b001110011101111 : data = 16'b0000000000111000;
            15'b001110011110000 : data = 16'b0000000000110111;
            15'b001110011110001 : data = 16'b0000000000110110;
            15'b001110011110010 : data = 16'b0000000000110101;
            15'b001110011110011 : data = 16'b0000000000110100;
            15'b001110011110100 : data = 16'b0000000000110011;
            15'b001110011110101 : data = 16'b0000000000110001;
            15'b001110011110110 : data = 16'b0000000000110000;
            15'b001110011110111 : data = 16'b0000000000101111;
            15'b001110011111000 : data = 16'b0000000000101110;
            15'b001110011111001 : data = 16'b0000000000101101;
            15'b001110011111010 : data = 16'b0000000000101100;
            15'b001110011111011 : data = 16'b0000000000101011;
            15'b001110011111100 : data = 16'b0000000000101010;
            15'b001110011111101 : data = 16'b0000000000101001;
            15'b001110011111110 : data = 16'b0000000000101000;
            15'b001110011111111 : data = 16'b0000000000100111;
            15'b001110100000000 : data = 16'b0000000000100110;
            15'b001110100000001 : data = 16'b0000000000100101;
            15'b001110100000010 : data = 16'b0000000000100100;
            15'b001110100000011 : data = 16'b0000000000100011;
            15'b001110100000100 : data = 16'b0000000000100010;
            15'b001110100000101 : data = 16'b0000000000100001;
            15'b001110100000110 : data = 16'b0000000000100000;
            15'b001110100000111 : data = 16'b0000000000011111;
            15'b001110100001000 : data = 16'b0000000000011110;
            15'b001110100001001 : data = 16'b0000000000011110;
            15'b001110100001010 : data = 16'b0000000000011101;
            15'b001110100001011 : data = 16'b0000000000011100;
            15'b001110100001100 : data = 16'b0000000000011011;
            15'b001110100001101 : data = 16'b0000000000011010;
            15'b001110100001110 : data = 16'b0000000000011001;
            15'b001110100001111 : data = 16'b0000000000011001;
            15'b001110100010000 : data = 16'b0000000000011000;
            15'b001110100010001 : data = 16'b0000000000010111;
            15'b001110100010010 : data = 16'b0000000000010110;
            15'b001110100010011 : data = 16'b0000000000010110;
            15'b001110100010100 : data = 16'b0000000000010101;
            15'b001110100010101 : data = 16'b0000000000010100;
            15'b001110100010110 : data = 16'b0000000000010011;
            15'b001110100010111 : data = 16'b0000000000010011;
            15'b001110100011000 : data = 16'b0000000000010010;
            15'b001110100011001 : data = 16'b0000000000010001;
            15'b001110100011010 : data = 16'b0000000000010001;
            15'b001110100011011 : data = 16'b0000000000010000;
            15'b001110100011100 : data = 16'b0000000000001111;
            15'b001110100011101 : data = 16'b0000000000001111;
            15'b001110100011110 : data = 16'b0000000000001110;
            15'b001110100011111 : data = 16'b0000000000001110;
            15'b001110100100000 : data = 16'b0000000000001101;
            15'b001110100100001 : data = 16'b0000000000001100;
            15'b001110100100010 : data = 16'b0000000000001100;
            15'b001110100100011 : data = 16'b0000000000001011;
            15'b001110100100100 : data = 16'b0000000000001011;
            15'b001110100100101 : data = 16'b0000000000001010;
            15'b001110100100110 : data = 16'b0000000000001010;
            15'b001110100100111 : data = 16'b0000000000001001;
            15'b001110100101000 : data = 16'b0000000000001001;
            15'b001110100101001 : data = 16'b0000000000001000;
            15'b001110100101010 : data = 16'b0000000000001000;
            15'b001110100101011 : data = 16'b0000000000001000;
            15'b001110100101100 : data = 16'b0000000000000111;
            15'b001110100101101 : data = 16'b0000000000000111;
            15'b001110100101110 : data = 16'b0000000000000110;
            15'b001110100101111 : data = 16'b0000000000000110;
            15'b001110100110000 : data = 16'b0000000000000110;
            15'b001110100110001 : data = 16'b0000000000000101;
            15'b001110100110010 : data = 16'b0000000000000101;
            15'b001110100110011 : data = 16'b0000000000000101;
            15'b001110100110100 : data = 16'b0000000000000100;
            15'b001110100110101 : data = 16'b0000000000000100;
            15'b001110100110110 : data = 16'b0000000000000100;
            15'b001110100110111 : data = 16'b0000000000000011;
            15'b001110100111000 : data = 16'b0000000000000011;
            15'b001110100111001 : data = 16'b0000000000000011;
            15'b001110100111010 : data = 16'b0000000000000011;
            15'b001110100111011 : data = 16'b0000000000000010;
            15'b001110100111100 : data = 16'b0000000000000010;
            15'b001110100111101 : data = 16'b0000000000000010;
            15'b001110100111110 : data = 16'b0000000000000010;
            15'b001110100111111 : data = 16'b0000000000000010;
            15'b001110101000000 : data = 16'b0000000000000001;
            15'b001110101000001 : data = 16'b0000000000000001;
            15'b001110101000010 : data = 16'b0000000000000001;
            15'b001110101000011 : data = 16'b0000000000000001;
            15'b001110101000100 : data = 16'b0000000000000001;
            15'b001110101000101 : data = 16'b0000000000000001;
            15'b001110101000110 : data = 16'b0000000000000001;
            15'b001110101000111 : data = 16'b0000000000000001;
            15'b001110101001000 : data = 16'b0000000000000001;
            15'b001110101001001 : data = 16'b0000000000000001;
            15'b001110101001010 : data = 16'b0000000000000001;
            15'b001110101001011 : data = 16'b0000000000000001;
            15'b001110101001100 : data = 16'b0000000000000001;
            15'b001110101001101 : data = 16'b0000000000000001;
            15'b001110101001110 : data = 16'b0000000000000001;
            15'b001110101001111 : data = 16'b0000000000000001;
            15'b001110101010000 : data = 16'b0000000000000001;
            15'b001110101010001 : data = 16'b0000000000000001;
            15'b001110101010010 : data = 16'b0000000000000001;
            15'b001110101010011 : data = 16'b0000000000000001;
            15'b001110101010100 : data = 16'b0000000000000001;
            15'b001110101010101 : data = 16'b0000000000000001;
            15'b001110101010110 : data = 16'b0000000000000001;
            15'b001110101010111 : data = 16'b0000000000000001;
            15'b001110101011000 : data = 16'b0000000000000001;
            15'b001110101011001 : data = 16'b0000000000000010;
            15'b001110101011010 : data = 16'b0000000000000010;
            15'b001110101011011 : data = 16'b0000000000000010;
            15'b001110101011100 : data = 16'b0000000000000010;
            15'b001110101011101 : data = 16'b0000000000000010;
            15'b001110101011110 : data = 16'b0000000000000011;
            15'b001110101011111 : data = 16'b0000000000000011;
            15'b001110101100000 : data = 16'b0000000000000011;
            15'b001110101100001 : data = 16'b0000000000000011;
            15'b001110101100010 : data = 16'b0000000000000100;
            15'b001110101100011 : data = 16'b0000000000000100;
            15'b001110101100100 : data = 16'b0000000000000100;
            15'b001110101100101 : data = 16'b0000000000000101;
            15'b001110101100110 : data = 16'b0000000000000101;
            15'b001110101100111 : data = 16'b0000000000000101;
            15'b001110101101000 : data = 16'b0000000000000110;
            15'b001110101101001 : data = 16'b0000000000000110;
            15'b001110101101010 : data = 16'b0000000000000110;
            15'b001110101101011 : data = 16'b0000000000000111;
            15'b001110101101100 : data = 16'b0000000000000111;
            15'b001110101101101 : data = 16'b0000000000001000;
            15'b001110101101110 : data = 16'b0000000000001000;
            15'b001110101101111 : data = 16'b0000000000001000;
            15'b001110101110000 : data = 16'b0000000000001001;
            15'b001110101110001 : data = 16'b0000000000001001;
            15'b001110101110010 : data = 16'b0000000000001010;
            15'b001110101110011 : data = 16'b0000000000001010;
            15'b001110101110100 : data = 16'b0000000000001011;
            15'b001110101110101 : data = 16'b0000000000001011;
            15'b001110101110110 : data = 16'b0000000000001100;
            15'b001110101110111 : data = 16'b0000000000001100;
            15'b001110101111000 : data = 16'b0000000000001101;
            15'b001110101111001 : data = 16'b0000000000001110;
            15'b001110101111010 : data = 16'b0000000000001110;
            15'b001110101111011 : data = 16'b0000000000001111;
            15'b001110101111100 : data = 16'b0000000000001111;
            15'b001110101111101 : data = 16'b0000000000010000;
            15'b001110101111110 : data = 16'b0000000000010001;
            15'b001110101111111 : data = 16'b0000000000010001;
            15'b001110110000000 : data = 16'b0000000000010010;
            15'b001110110000001 : data = 16'b0000000000010011;
            15'b001110110000010 : data = 16'b0000000000010011;
            15'b001110110000011 : data = 16'b0000000000010100;
            15'b001110110000100 : data = 16'b0000000000010101;
            15'b001110110000101 : data = 16'b0000000000010110;
            15'b001110110000110 : data = 16'b0000000000010110;
            15'b001110110000111 : data = 16'b0000000000010111;
            15'b001110110001000 : data = 16'b0000000000011000;
            15'b001110110001001 : data = 16'b0000000000011001;
            15'b001110110001010 : data = 16'b0000000000011001;
            15'b001110110001011 : data = 16'b0000000000011010;
            15'b001110110001100 : data = 16'b0000000000011011;
            15'b001110110001101 : data = 16'b0000000000011100;
            15'b001110110001110 : data = 16'b0000000000011101;
            15'b001110110001111 : data = 16'b0000000000011110;
            15'b001110110010000 : data = 16'b0000000000011110;
            15'b001110110010001 : data = 16'b0000000000011111;
            15'b001110110010010 : data = 16'b0000000000100000;
            15'b001110110010011 : data = 16'b0000000000100001;
            15'b001110110010100 : data = 16'b0000000000100010;
            15'b001110110010101 : data = 16'b0000000000100011;
            15'b001110110010110 : data = 16'b0000000000100100;
            15'b001110110010111 : data = 16'b0000000000100101;
            15'b001110110011000 : data = 16'b0000000000100110;
            15'b001110110011001 : data = 16'b0000000000100111;
            15'b001110110011010 : data = 16'b0000000000101000;
            15'b001110110011011 : data = 16'b0000000000101001;
            15'b001110110011100 : data = 16'b0000000000101010;
            15'b001110110011101 : data = 16'b0000000000101011;
            15'b001110110011110 : data = 16'b0000000000101100;
            15'b001110110011111 : data = 16'b0000000000101101;
            15'b001110110100000 : data = 16'b0000000000101110;
            15'b001110110100001 : data = 16'b0000000000101111;
            15'b001110110100010 : data = 16'b0000000000110000;
            15'b001110110100011 : data = 16'b0000000000110001;
            15'b001110110100100 : data = 16'b0000000000110011;
            15'b001110110100101 : data = 16'b0000000000110100;
            15'b001110110100110 : data = 16'b0000000000110101;
            15'b001110110100111 : data = 16'b0000000000110110;
            15'b001110110101000 : data = 16'b0000000000110111;
            15'b001110110101001 : data = 16'b0000000000111000;
            15'b001110110101010 : data = 16'b0000000000111010;
            15'b001110110101011 : data = 16'b0000000000111011;
            15'b001110110101100 : data = 16'b0000000000111100;
            15'b001110110101101 : data = 16'b0000000000111101;
            15'b001110110101110 : data = 16'b0000000000111111;
            15'b001110110101111 : data = 16'b0000000001000000;
            15'b001110110110000 : data = 16'b0000000001000001;
            15'b001110110110001 : data = 16'b0000000001000010;
            15'b001110110110010 : data = 16'b0000000001000100;
            15'b001110110110011 : data = 16'b0000000001000101;
            15'b001110110110100 : data = 16'b0000000001000110;
            15'b001110110110101 : data = 16'b0000000001001000;
            15'b001110110110110 : data = 16'b0000000001001001;
            15'b001110110110111 : data = 16'b0000000001001011;
            15'b001110110111000 : data = 16'b0000000001001100;
            15'b001110110111001 : data = 16'b0000000001001101;
            15'b001110110111010 : data = 16'b0000000001001111;
            15'b001110110111011 : data = 16'b0000000001010000;
            15'b001110110111100 : data = 16'b0000000001010010;
            15'b001110110111101 : data = 16'b0000000001010011;
            15'b001110110111110 : data = 16'b0000000001010101;
            15'b001110110111111 : data = 16'b0000000001010110;
            15'b001110111000000 : data = 16'b0000000001010111;
            15'b001110111000001 : data = 16'b0000000001011001;
            15'b001110111000010 : data = 16'b0000000001011011;
            15'b001110111000011 : data = 16'b0000000001011100;
            15'b001110111000100 : data = 16'b0000000001011110;
            15'b001110111000101 : data = 16'b0000000001011111;
            15'b001110111000110 : data = 16'b0000000001100001;
            15'b001110111000111 : data = 16'b0000000001100010;
            15'b001110111001000 : data = 16'b0000000001100100;
            15'b001110111001001 : data = 16'b0000000001100110;
            15'b001110111001010 : data = 16'b0000000001100111;
            15'b001110111001011 : data = 16'b0000000001101001;
            15'b001110111001100 : data = 16'b0000000001101010;
            15'b001110111001101 : data = 16'b0000000001101100;
            15'b001110111001110 : data = 16'b0000000001101110;
            15'b001110111001111 : data = 16'b0000000001101111;
            15'b001110111010000 : data = 16'b0000000001110001;
            15'b001110111010001 : data = 16'b0000000001110011;
            15'b001110111010010 : data = 16'b0000000001110101;
            15'b001110111010011 : data = 16'b0000000001110110;
            15'b001110111010100 : data = 16'b0000000001111000;
            15'b001110111010101 : data = 16'b0000000001111010;
            15'b001110111010110 : data = 16'b0000000001111100;
            15'b001110111010111 : data = 16'b0000000001111101;
            15'b001110111011000 : data = 16'b0000000001111111;
            15'b001110111011001 : data = 16'b0000000010000001;
            15'b001110111011010 : data = 16'b0000000010000011;
            15'b001110111011011 : data = 16'b0000000010000101;
            15'b001110111011100 : data = 16'b0000000010000111;
            15'b001110111011101 : data = 16'b0000000010001000;
            15'b001110111011110 : data = 16'b0000000010001010;
            15'b001110111011111 : data = 16'b0000000010001100;
            15'b001110111100000 : data = 16'b0000000010001110;
            15'b001110111100001 : data = 16'b0000000010010000;
            15'b001110111100010 : data = 16'b0000000010010010;
            15'b001110111100011 : data = 16'b0000000010010100;
            15'b001110111100100 : data = 16'b0000000010010110;
            15'b001110111100101 : data = 16'b0000000010011000;
            15'b001110111100110 : data = 16'b0000000010011010;
            15'b001110111100111 : data = 16'b0000000010011100;
            15'b001110111101000 : data = 16'b0000000010011110;
            15'b001110111101001 : data = 16'b0000000010100000;
            15'b001110111101010 : data = 16'b0000000010100010;
            15'b001110111101011 : data = 16'b0000000010100100;
            15'b001110111101100 : data = 16'b0000000010100110;
            15'b001110111101101 : data = 16'b0000000010101000;
            15'b001110111101110 : data = 16'b0000000010101010;
            15'b001110111101111 : data = 16'b0000000010101100;
            15'b001110111110000 : data = 16'b0000000010101110;
            15'b001110111110001 : data = 16'b0000000010110000;
            15'b001110111110010 : data = 16'b0000000010110011;
            15'b001110111110011 : data = 16'b0000000010110101;
            15'b001110111110100 : data = 16'b0000000010110111;
            15'b001110111110101 : data = 16'b0000000010111001;
            15'b001110111110110 : data = 16'b0000000010111011;
            15'b001110111110111 : data = 16'b0000000010111101;
            15'b001110111111000 : data = 16'b0000000011000000;
            15'b001110111111001 : data = 16'b0000000011000010;
            15'b001110111111010 : data = 16'b0000000011000100;
            15'b001110111111011 : data = 16'b0000000011000110;
            15'b001110111111100 : data = 16'b0000000011001001;
            15'b001110111111101 : data = 16'b0000000011001011;
            15'b001110111111110 : data = 16'b0000000011001101;
            15'b001110111111111 : data = 16'b0000000011010000;
            15'b001111000000000 : data = 16'b0000000011010010;
            15'b001111000000001 : data = 16'b0000000011010100;
            15'b001111000000010 : data = 16'b0000000011010111;
            15'b001111000000011 : data = 16'b0000000011011001;
            15'b001111000000100 : data = 16'b0000000011011011;
            15'b001111000000101 : data = 16'b0000000011011110;
            15'b001111000000110 : data = 16'b0000000011100000;
            15'b001111000000111 : data = 16'b0000000011100010;
            15'b001111000001000 : data = 16'b0000000011100101;
            15'b001111000001001 : data = 16'b0000000011100111;
            15'b001111000001010 : data = 16'b0000000011101010;
            15'b001111000001011 : data = 16'b0000000011101100;
            15'b001111000001100 : data = 16'b0000000011101111;
            15'b001111000001101 : data = 16'b0000000011110001;
            15'b001111000001110 : data = 16'b0000000011110100;
            15'b001111000001111 : data = 16'b0000000011110110;
            15'b001111000010000 : data = 16'b0000000011111001;
            15'b001111000010001 : data = 16'b0000000011111011;
            15'b001111000010010 : data = 16'b0000000011111110;
            15'b001111000010011 : data = 16'b0000000100000000;
            15'b001111000010100 : data = 16'b0000000100000011;
            15'b001111000010101 : data = 16'b0000000100000101;
            15'b001111000010110 : data = 16'b0000000100001000;
            15'b001111000010111 : data = 16'b0000000100001011;
            15'b001111000011000 : data = 16'b0000000100001101;
            15'b001111000011001 : data = 16'b0000000100010000;
            15'b001111000011010 : data = 16'b0000000100010011;
            15'b001111000011011 : data = 16'b0000000100010101;
            15'b001111000011100 : data = 16'b0000000100011000;
            15'b001111000011101 : data = 16'b0000000100011011;
            15'b001111000011110 : data = 16'b0000000100011101;
            15'b001111000011111 : data = 16'b0000000100100000;
            15'b001111000100000 : data = 16'b0000000100100011;
            15'b001111000100001 : data = 16'b0000000100100110;
            15'b001111000100010 : data = 16'b0000000100101000;
            15'b001111000100011 : data = 16'b0000000100101011;
            15'b001111000100100 : data = 16'b0000000100101110;
            15'b001111000100101 : data = 16'b0000000100110001;
            15'b001111000100110 : data = 16'b0000000100110011;
            15'b001111000100111 : data = 16'b0000000100110110;
            15'b001111000101000 : data = 16'b0000000100111001;
            15'b001111000101001 : data = 16'b0000000100111100;
            15'b001111000101010 : data = 16'b0000000100111111;
            15'b001111000101011 : data = 16'b0000000101000010;
            15'b001111000101100 : data = 16'b0000000101000101;
            15'b001111000101101 : data = 16'b0000000101000111;
            15'b001111000101110 : data = 16'b0000000101001010;
            15'b001111000101111 : data = 16'b0000000101001101;
            15'b001111000110000 : data = 16'b0000000101010000;
            15'b001111000110001 : data = 16'b0000000101010011;
            15'b001111000110010 : data = 16'b0000000101010110;
            15'b001111000110011 : data = 16'b0000000101011001;
            15'b001111000110100 : data = 16'b0000000101011100;
            15'b001111000110101 : data = 16'b0000000101011111;
            15'b001111000110110 : data = 16'b0000000101100010;
            15'b001111000110111 : data = 16'b0000000101100101;
            15'b001111000111000 : data = 16'b0000000101101000;
            15'b001111000111001 : data = 16'b0000000101101011;
            15'b001111000111010 : data = 16'b0000000101101110;
            15'b001111000111011 : data = 16'b0000000101110001;
            15'b001111000111100 : data = 16'b0000000101110100;
            15'b001111000111101 : data = 16'b0000000101110111;
            15'b001111000111110 : data = 16'b0000000101111011;
            15'b001111000111111 : data = 16'b0000000101111110;
            15'b001111001000000 : data = 16'b0000000110000001;
            15'b001111001000001 : data = 16'b0000000110000100;
            15'b001111001000010 : data = 16'b0000000110000111;
            15'b001111001000011 : data = 16'b0000000110001010;
            15'b001111001000100 : data = 16'b0000000110001110;
            15'b001111001000101 : data = 16'b0000000110010001;
            15'b001111001000110 : data = 16'b0000000110010100;
            15'b001111001000111 : data = 16'b0000000110010111;
            15'b001111001001000 : data = 16'b0000000110011010;
            15'b001111001001001 : data = 16'b0000000110011110;
            15'b001111001001010 : data = 16'b0000000110100001;
            15'b001111001001011 : data = 16'b0000000110100100;
            15'b001111001001100 : data = 16'b0000000110100111;
            15'b001111001001101 : data = 16'b0000000110101011;
            15'b001111001001110 : data = 16'b0000000110101110;
            15'b001111001001111 : data = 16'b0000000110110001;
            15'b001111001010000 : data = 16'b0000000110110101;
            15'b001111001010001 : data = 16'b0000000110111000;
            15'b001111001010010 : data = 16'b0000000110111011;
            15'b001111001010011 : data = 16'b0000000110111111;
            15'b001111001010100 : data = 16'b0000000111000010;
            15'b001111001010101 : data = 16'b0000000111000110;
            15'b001111001010110 : data = 16'b0000000111001001;
            15'b001111001010111 : data = 16'b0000000111001101;
            15'b001111001011000 : data = 16'b0000000111010000;
            15'b001111001011001 : data = 16'b0000000111010011;
            15'b001111001011010 : data = 16'b0000000111010111;
            15'b001111001011011 : data = 16'b0000000111011010;
            15'b001111001011100 : data = 16'b0000000111011110;
            15'b001111001011101 : data = 16'b0000000111100001;
            15'b001111001011110 : data = 16'b0000000111100101;
            15'b001111001011111 : data = 16'b0000000111101000;
            15'b001111001100000 : data = 16'b0000000111101100;
            15'b001111001100001 : data = 16'b0000000111110000;
            15'b001111001100010 : data = 16'b0000000111110011;
            15'b001111001100011 : data = 16'b0000000111110111;
            15'b001111001100100 : data = 16'b0000000111111010;
            15'b001111001100101 : data = 16'b0000000111111110;
            15'b001111001100110 : data = 16'b0000001000000010;
            15'b001111001100111 : data = 16'b0000001000000101;
            15'b001111001101000 : data = 16'b0000001000001001;
            15'b001111001101001 : data = 16'b0000001000001100;
            15'b001111001101010 : data = 16'b0000001000010000;
            15'b001111001101011 : data = 16'b0000001000010100;
            15'b001111001101100 : data = 16'b0000001000011000;
            15'b001111001101101 : data = 16'b0000001000011011;
            15'b001111001101110 : data = 16'b0000001000011111;
            15'b001111001101111 : data = 16'b0000001000100011;
            15'b001111001110000 : data = 16'b0000001000100110;
            15'b001111001110001 : data = 16'b0000001000101010;
            15'b001111001110010 : data = 16'b0000001000101110;
            15'b001111001110011 : data = 16'b0000001000110010;
            15'b001111001110100 : data = 16'b0000001000110110;
            15'b001111001110101 : data = 16'b0000001000111001;
            15'b001111001110110 : data = 16'b0000001000111101;
            15'b001111001110111 : data = 16'b0000001001000001;
            15'b001111001111000 : data = 16'b0000001001000101;
            15'b001111001111001 : data = 16'b0000001001001001;
            15'b001111001111010 : data = 16'b0000001001001101;
            15'b001111001111011 : data = 16'b0000001001010001;
            15'b001111001111100 : data = 16'b0000001001010100;
            15'b001111001111101 : data = 16'b0000001001011000;
            15'b001111001111110 : data = 16'b0000001001011100;
            15'b001111001111111 : data = 16'b0000001001100000;
            15'b001111010000000 : data = 16'b0000001001100100;
            15'b001111010000001 : data = 16'b0000001001101000;
            15'b001111010000010 : data = 16'b0000001001101100;
            15'b001111010000011 : data = 16'b0000001001110000;
            15'b001111010000100 : data = 16'b0000001001110100;
            15'b001111010000101 : data = 16'b0000001001111000;
            15'b001111010000110 : data = 16'b0000001001111100;
            15'b001111010000111 : data = 16'b0000001010000000;
            15'b001111010001000 : data = 16'b0000001010000100;
            15'b001111010001001 : data = 16'b0000001010001000;
            15'b001111010001010 : data = 16'b0000001010001100;
            15'b001111010001011 : data = 16'b0000001010010000;
            15'b001111010001100 : data = 16'b0000001010010101;
            15'b001111010001101 : data = 16'b0000001010011001;
            15'b001111010001110 : data = 16'b0000001010011101;
            15'b001111010001111 : data = 16'b0000001010100001;
            15'b001111010010000 : data = 16'b0000001010100101;
            15'b001111010010001 : data = 16'b0000001010101001;
            15'b001111010010010 : data = 16'b0000001010101101;
            15'b001111010010011 : data = 16'b0000001010110010;
            15'b001111010010100 : data = 16'b0000001010110110;
            15'b001111010010101 : data = 16'b0000001010111010;
            15'b001111010010110 : data = 16'b0000001010111110;
            15'b001111010010111 : data = 16'b0000001011000011;
            15'b001111010011000 : data = 16'b0000001011000111;
            15'b001111010011001 : data = 16'b0000001011001011;
            15'b001111010011010 : data = 16'b0000001011001111;
            15'b001111010011011 : data = 16'b0000001011010100;
            15'b001111010011100 : data = 16'b0000001011011000;
            15'b001111010011101 : data = 16'b0000001011011100;
            15'b001111010011110 : data = 16'b0000001011100001;
            15'b001111010011111 : data = 16'b0000001011100101;
            15'b001111010100000 : data = 16'b0000001011101001;
            15'b001111010100001 : data = 16'b0000001011101110;
            15'b001111010100010 : data = 16'b0000001011110010;
            15'b001111010100011 : data = 16'b0000001011110111;
            15'b001111010100100 : data = 16'b0000001011111011;
            15'b001111010100101 : data = 16'b0000001011111111;
            15'b001111010100110 : data = 16'b0000001100000100;
            15'b001111010100111 : data = 16'b0000001100001000;
            15'b001111010101000 : data = 16'b0000001100001101;
            15'b001111010101001 : data = 16'b0000001100010001;
            15'b001111010101010 : data = 16'b0000001100010110;
            15'b001111010101011 : data = 16'b0000001100011010;
            15'b001111010101100 : data = 16'b0000001100011111;
            15'b001111010101101 : data = 16'b0000001100100011;
            15'b001111010101110 : data = 16'b0000001100101000;
            15'b001111010101111 : data = 16'b0000001100101100;
            15'b001111010110000 : data = 16'b0000001100110001;
            15'b001111010110001 : data = 16'b0000001100110101;
            15'b001111010110010 : data = 16'b0000001100111010;
            15'b001111010110011 : data = 16'b0000001100111111;
            15'b001111010110100 : data = 16'b0000001101000011;
            15'b001111010110101 : data = 16'b0000001101001000;
            15'b001111010110110 : data = 16'b0000001101001100;
            15'b001111010110111 : data = 16'b0000001101010001;
            15'b001111010111000 : data = 16'b0000001101010110;
            15'b001111010111001 : data = 16'b0000001101011010;
            15'b001111010111010 : data = 16'b0000001101011111;
            15'b001111010111011 : data = 16'b0000001101100100;
            15'b001111010111100 : data = 16'b0000001101101001;
            15'b001111010111101 : data = 16'b0000001101101101;
            15'b001111010111110 : data = 16'b0000001101110010;
            15'b001111010111111 : data = 16'b0000001101110111;
            15'b001111011000000 : data = 16'b0000001101111011;
            15'b001111011000001 : data = 16'b0000001110000000;
            15'b001111011000010 : data = 16'b0000001110000101;
            15'b001111011000011 : data = 16'b0000001110001010;
            15'b001111011000100 : data = 16'b0000001110001111;
            15'b001111011000101 : data = 16'b0000001110010011;
            15'b001111011000110 : data = 16'b0000001110011000;
            15'b001111011000111 : data = 16'b0000001110011101;
            15'b001111011001000 : data = 16'b0000001110100010;
            15'b001111011001001 : data = 16'b0000001110100111;
            15'b001111011001010 : data = 16'b0000001110101100;
            15'b001111011001011 : data = 16'b0000001110110001;
            15'b001111011001100 : data = 16'b0000001110110110;
            15'b001111011001101 : data = 16'b0000001110111011;
            15'b001111011001110 : data = 16'b0000001110111111;
            15'b001111011001111 : data = 16'b0000001111000100;
            15'b001111011010000 : data = 16'b0000001111001001;
            15'b001111011010001 : data = 16'b0000001111001110;
            15'b001111011010010 : data = 16'b0000001111010011;
            15'b001111011010011 : data = 16'b0000001111011000;
            15'b001111011010100 : data = 16'b0000001111011101;
            15'b001111011010101 : data = 16'b0000001111100010;
            15'b001111011010110 : data = 16'b0000001111100111;
            15'b001111011010111 : data = 16'b0000001111101100;
            15'b001111011011000 : data = 16'b0000001111110010;
            15'b001111011011001 : data = 16'b0000001111110111;
            15'b001111011011010 : data = 16'b0000001111111100;
            15'b001111011011011 : data = 16'b0000010000000001;
            15'b001111011011100 : data = 16'b0000010000000110;
            15'b001111011011101 : data = 16'b0000010000001011;
            15'b001111011011110 : data = 16'b0000010000010000;
            15'b001111011011111 : data = 16'b0000010000010101;
            15'b001111011100000 : data = 16'b0000010000011011;
            15'b001111011100001 : data = 16'b0000010000100000;
            15'b001111011100010 : data = 16'b0000010000100101;
            15'b001111011100011 : data = 16'b0000010000101010;
            15'b001111011100100 : data = 16'b0000010000101111;
            15'b001111011100101 : data = 16'b0000010000110101;
            15'b001111011100110 : data = 16'b0000010000111010;
            15'b001111011100111 : data = 16'b0000010000111111;
            15'b001111011101000 : data = 16'b0000010001000100;
            15'b001111011101001 : data = 16'b0000010001001010;
            15'b001111011101010 : data = 16'b0000010001001111;
            15'b001111011101011 : data = 16'b0000010001010100;
            15'b001111011101100 : data = 16'b0000010001011001;
            15'b001111011101101 : data = 16'b0000010001011111;
            15'b001111011101110 : data = 16'b0000010001100100;
            15'b001111011101111 : data = 16'b0000010001101001;
            15'b001111011110000 : data = 16'b0000010001101111;
            15'b001111011110001 : data = 16'b0000010001110100;
            15'b001111011110010 : data = 16'b0000010001111010;
            15'b001111011110011 : data = 16'b0000010001111111;
            15'b001111011110100 : data = 16'b0000010010000100;
            15'b001111011110101 : data = 16'b0000010010001010;
            15'b001111011110110 : data = 16'b0000010010001111;
            15'b001111011110111 : data = 16'b0000010010010101;
            15'b001111011111000 : data = 16'b0000010010011010;
            15'b001111011111001 : data = 16'b0000010010100000;
            15'b001111011111010 : data = 16'b0000010010100101;
            15'b001111011111011 : data = 16'b0000010010101011;
            15'b001111011111100 : data = 16'b0000010010110000;
            15'b001111011111101 : data = 16'b0000010010110110;
            15'b001111011111110 : data = 16'b0000010010111011;
            15'b001111011111111 : data = 16'b0000010011000001;
            15'b001111100000000 : data = 16'b0000010011000110;
            15'b001111100000001 : data = 16'b0000010011001100;
            15'b001111100000010 : data = 16'b0000010011010010;
            15'b001111100000011 : data = 16'b0000010011010111;
            15'b001111100000100 : data = 16'b0000010011011101;
            15'b001111100000101 : data = 16'b0000010011100010;
            15'b001111100000110 : data = 16'b0000010011101000;
            15'b001111100000111 : data = 16'b0000010011101110;
            15'b001111100001000 : data = 16'b0000010011110011;
            15'b001111100001001 : data = 16'b0000010011111001;
            15'b001111100001010 : data = 16'b0000010011111111;
            15'b001111100001011 : data = 16'b0000010100000100;
            15'b001111100001100 : data = 16'b0000010100001010;
            15'b001111100001101 : data = 16'b0000010100010000;
            15'b001111100001110 : data = 16'b0000010100010110;
            15'b001111100001111 : data = 16'b0000010100011011;
            15'b001111100010000 : data = 16'b0000010100100001;
            15'b001111100010001 : data = 16'b0000010100100111;
            15'b001111100010010 : data = 16'b0000010100101101;
            15'b001111100010011 : data = 16'b0000010100110010;
            15'b001111100010100 : data = 16'b0000010100111000;
            15'b001111100010101 : data = 16'b0000010100111110;
            15'b001111100010110 : data = 16'b0000010101000100;
            15'b001111100010111 : data = 16'b0000010101001010;
            15'b001111100011000 : data = 16'b0000010101010000;
            15'b001111100011001 : data = 16'b0000010101010101;
            15'b001111100011010 : data = 16'b0000010101011011;
            15'b001111100011011 : data = 16'b0000010101100001;
            15'b001111100011100 : data = 16'b0000010101100111;
            15'b001111100011101 : data = 16'b0000010101101101;
            15'b001111100011110 : data = 16'b0000010101110011;
            15'b001111100011111 : data = 16'b0000010101111001;
            15'b001111100100000 : data = 16'b0000010101111111;
            15'b001111100100001 : data = 16'b0000010110000101;
            15'b001111100100010 : data = 16'b0000010110001011;
            15'b001111100100011 : data = 16'b0000010110010001;
            15'b001111100100100 : data = 16'b0000010110010111;
            15'b001111100100101 : data = 16'b0000010110011101;
            15'b001111100100110 : data = 16'b0000010110100011;
            15'b001111100100111 : data = 16'b0000010110101001;
            15'b001111100101000 : data = 16'b0000010110101111;
            15'b001111100101001 : data = 16'b0000010110110101;
            15'b001111100101010 : data = 16'b0000010110111011;
            15'b001111100101011 : data = 16'b0000010111000001;
            15'b001111100101100 : data = 16'b0000010111000111;
            15'b001111100101101 : data = 16'b0000010111001110;
            15'b001111100101110 : data = 16'b0000010111010100;
            15'b001111100101111 : data = 16'b0000010111011010;
            15'b001111100110000 : data = 16'b0000010111100000;
            15'b001111100110001 : data = 16'b0000010111100110;
            15'b001111100110010 : data = 16'b0000010111101100;
            15'b001111100110011 : data = 16'b0000010111110011;
            15'b001111100110100 : data = 16'b0000010111111001;
            15'b001111100110101 : data = 16'b0000010111111111;
            15'b001111100110110 : data = 16'b0000011000000101;
            15'b001111100110111 : data = 16'b0000011000001011;
            15'b001111100111000 : data = 16'b0000011000010010;
            15'b001111100111001 : data = 16'b0000011000011000;
            15'b001111100111010 : data = 16'b0000011000011110;
            15'b001111100111011 : data = 16'b0000011000100101;
            15'b001111100111100 : data = 16'b0000011000101011;
            15'b001111100111101 : data = 16'b0000011000110001;
            15'b001111100111110 : data = 16'b0000011000111000;
            15'b001111100111111 : data = 16'b0000011000111110;
            15'b001111101000000 : data = 16'b0000011001000100;
            15'b001111101000001 : data = 16'b0000011001001011;
            15'b001111101000010 : data = 16'b0000011001010001;
            15'b001111101000011 : data = 16'b0000011001010111;
            15'b001111101000100 : data = 16'b0000011001011110;
            15'b001111101000101 : data = 16'b0000011001100100;
            15'b001111101000110 : data = 16'b0000011001101011;
            15'b001111101000111 : data = 16'b0000011001110001;
            15'b001111101001000 : data = 16'b0000011001111000;
            15'b001111101001001 : data = 16'b0000011001111110;
            15'b001111101001010 : data = 16'b0000011010000100;
            15'b001111101001011 : data = 16'b0000011010001011;
            15'b001111101001100 : data = 16'b0000011010010001;
            15'b001111101001101 : data = 16'b0000011010011000;
            15'b001111101001110 : data = 16'b0000011010011111;
            15'b001111101001111 : data = 16'b0000011010100101;
            15'b001111101010000 : data = 16'b0000011010101100;
            15'b001111101010001 : data = 16'b0000011010110010;
            15'b001111101010010 : data = 16'b0000011010111001;
            15'b001111101010011 : data = 16'b0000011010111111;
            15'b001111101010100 : data = 16'b0000011011000110;
            15'b001111101010101 : data = 16'b0000011011001101;
            15'b001111101010110 : data = 16'b0000011011010011;
            15'b001111101010111 : data = 16'b0000011011011010;
            15'b001111101011000 : data = 16'b0000011011100000;
            15'b001111101011001 : data = 16'b0000011011100111;
            15'b001111101011010 : data = 16'b0000011011101110;
            15'b001111101011011 : data = 16'b0000011011110100;
            15'b001111101011100 : data = 16'b0000011011111011;
            15'b001111101011101 : data = 16'b0000011100000010;
            15'b001111101011110 : data = 16'b0000011100001001;
            15'b001111101011111 : data = 16'b0000011100001111;
            15'b001111101100000 : data = 16'b0000011100010110;
            15'b001111101100001 : data = 16'b0000011100011101;
            15'b001111101100010 : data = 16'b0000011100100100;
            15'b001111101100011 : data = 16'b0000011100101010;
            15'b001111101100100 : data = 16'b0000011100110001;
            15'b001111101100101 : data = 16'b0000011100111000;
            15'b001111101100110 : data = 16'b0000011100111111;
            15'b001111101100111 : data = 16'b0000011101000110;
            15'b001111101101000 : data = 16'b0000011101001101;
            15'b001111101101001 : data = 16'b0000011101010011;
            15'b001111101101010 : data = 16'b0000011101011010;
            15'b001111101101011 : data = 16'b0000011101100001;
            15'b001111101101100 : data = 16'b0000011101101000;
            15'b001111101101101 : data = 16'b0000011101101111;
            15'b001111101101110 : data = 16'b0000011101110110;
            15'b001111101101111 : data = 16'b0000011101111101;
            15'b001111101110000 : data = 16'b0000011110000100;
            15'b001111101110001 : data = 16'b0000011110001011;
            15'b001111101110010 : data = 16'b0000011110010010;
            15'b001111101110011 : data = 16'b0000011110011001;
            15'b001111101110100 : data = 16'b0000011110100000;
            15'b001111101110101 : data = 16'b0000011110100111;
            15'b001111101110110 : data = 16'b0000011110101110;
            15'b001111101110111 : data = 16'b0000011110110101;
            15'b001111101111000 : data = 16'b0000011110111100;
            15'b001111101111001 : data = 16'b0000011111000011;
            15'b001111101111010 : data = 16'b0000011111001010;
            15'b001111101111011 : data = 16'b0000011111010001;
            15'b001111101111100 : data = 16'b0000011111011000;
            15'b001111101111101 : data = 16'b0000011111011111;
            15'b001111101111110 : data = 16'b0000011111100110;
            15'b001111101111111 : data = 16'b0000011111101101;
            15'b001111110000000 : data = 16'b0000011111110100;
            15'b001111110000001 : data = 16'b0000011111111100;
            15'b001111110000010 : data = 16'b0000100000000011;
            15'b001111110000011 : data = 16'b0000100000001010;
            15'b001111110000100 : data = 16'b0000100000010001;
            15'b001111110000101 : data = 16'b0000100000011000;
            15'b001111110000110 : data = 16'b0000100000100000;
            15'b001111110000111 : data = 16'b0000100000100111;
            15'b001111110001000 : data = 16'b0000100000101110;
            15'b001111110001001 : data = 16'b0000100000110101;
            15'b001111110001010 : data = 16'b0000100000111101;
            15'b001111110001011 : data = 16'b0000100001000100;
            15'b001111110001100 : data = 16'b0000100001001011;
            15'b001111110001101 : data = 16'b0000100001010010;
            15'b001111110001110 : data = 16'b0000100001011010;
            15'b001111110001111 : data = 16'b0000100001100001;
            15'b001111110010000 : data = 16'b0000100001101000;
            15'b001111110010001 : data = 16'b0000100001110000;
            15'b001111110010010 : data = 16'b0000100001110111;
            15'b001111110010011 : data = 16'b0000100001111110;
            15'b001111110010100 : data = 16'b0000100010000110;
            15'b001111110010101 : data = 16'b0000100010001101;
            15'b001111110010110 : data = 16'b0000100010010101;
            15'b001111110010111 : data = 16'b0000100010011100;
            15'b001111110011000 : data = 16'b0000100010100011;
            15'b001111110011001 : data = 16'b0000100010101011;
            15'b001111110011010 : data = 16'b0000100010110010;
            15'b001111110011011 : data = 16'b0000100010111010;
            15'b001111110011100 : data = 16'b0000100011000001;
            15'b001111110011101 : data = 16'b0000100011001001;
            15'b001111110011110 : data = 16'b0000100011010000;
            15'b001111110011111 : data = 16'b0000100011011000;
            15'b001111110100000 : data = 16'b0000100011011111;
            15'b001111110100001 : data = 16'b0000100011100111;
            15'b001111110100010 : data = 16'b0000100011101110;
            15'b001111110100011 : data = 16'b0000100011110110;
            15'b001111110100100 : data = 16'b0000100011111110;
            15'b001111110100101 : data = 16'b0000100100000101;
            15'b001111110100110 : data = 16'b0000100100001101;
            15'b001111110100111 : data = 16'b0000100100010100;
            15'b001111110101000 : data = 16'b0000100100011100;
            15'b001111110101001 : data = 16'b0000100100100100;
            15'b001111110101010 : data = 16'b0000100100101011;
            15'b001111110101011 : data = 16'b0000100100110011;
            15'b001111110101100 : data = 16'b0000100100111011;
            15'b001111110101101 : data = 16'b0000100101000010;
            15'b001111110101110 : data = 16'b0000100101001010;
            15'b001111110101111 : data = 16'b0000100101010010;
            15'b001111110110000 : data = 16'b0000100101011001;
            15'b001111110110001 : data = 16'b0000100101100001;
            15'b001111110110010 : data = 16'b0000100101101001;
            15'b001111110110011 : data = 16'b0000100101110001;
            15'b001111110110100 : data = 16'b0000100101111000;
            15'b001111110110101 : data = 16'b0000100110000000;
            15'b001111110110110 : data = 16'b0000100110001000;
            15'b001111110110111 : data = 16'b0000100110010000;
            15'b001111110111000 : data = 16'b0000100110010111;
            15'b001111110111001 : data = 16'b0000100110011111;
            15'b001111110111010 : data = 16'b0000100110100111;
            15'b001111110111011 : data = 16'b0000100110101111;
            15'b001111110111100 : data = 16'b0000100110110111;
            15'b001111110111101 : data = 16'b0000100110111111;
            15'b001111110111110 : data = 16'b0000100111000111;
            15'b001111110111111 : data = 16'b0000100111001111;
            15'b001111111000000 : data = 16'b0000100111010110;
            15'b001111111000001 : data = 16'b0000100111011110;
            15'b001111111000010 : data = 16'b0000100111100110;
            15'b001111111000011 : data = 16'b0000100111101110;
            15'b001111111000100 : data = 16'b0000100111110110;
            15'b001111111000101 : data = 16'b0000100111111110;
            15'b001111111000110 : data = 16'b0000101000000110;
            15'b001111111000111 : data = 16'b0000101000001110;
            15'b001111111001000 : data = 16'b0000101000010110;
            15'b001111111001001 : data = 16'b0000101000011110;
            15'b001111111001010 : data = 16'b0000101000100110;
            15'b001111111001011 : data = 16'b0000101000101110;
            15'b001111111001100 : data = 16'b0000101000110110;
            15'b001111111001101 : data = 16'b0000101000111110;
            15'b001111111001110 : data = 16'b0000101001000110;
            15'b001111111001111 : data = 16'b0000101001001110;
            15'b001111111010000 : data = 16'b0000101001010111;
            15'b001111111010001 : data = 16'b0000101001011111;
            15'b001111111010010 : data = 16'b0000101001100111;
            15'b001111111010011 : data = 16'b0000101001101111;
            15'b001111111010100 : data = 16'b0000101001110111;
            15'b001111111010101 : data = 16'b0000101001111111;
            15'b001111111010110 : data = 16'b0000101010000111;
            15'b001111111010111 : data = 16'b0000101010010000;
            15'b001111111011000 : data = 16'b0000101010011000;
            15'b001111111011001 : data = 16'b0000101010100000;
            15'b001111111011010 : data = 16'b0000101010101000;
            15'b001111111011011 : data = 16'b0000101010110000;
            15'b001111111011100 : data = 16'b0000101010111001;
            15'b001111111011101 : data = 16'b0000101011000001;
            15'b001111111011110 : data = 16'b0000101011001001;
            15'b001111111011111 : data = 16'b0000101011010010;
            15'b001111111100000 : data = 16'b0000101011011010;
            15'b001111111100001 : data = 16'b0000101011100010;
            15'b001111111100010 : data = 16'b0000101011101010;
            15'b001111111100011 : data = 16'b0000101011110011;
            15'b001111111100100 : data = 16'b0000101011111011;
            15'b001111111100101 : data = 16'b0000101100000011;
            15'b001111111100110 : data = 16'b0000101100001100;
            15'b001111111100111 : data = 16'b0000101100010100;
            15'b001111111101000 : data = 16'b0000101100011101;
            15'b001111111101001 : data = 16'b0000101100100101;
            15'b001111111101010 : data = 16'b0000101100101101;
            15'b001111111101011 : data = 16'b0000101100110110;
            15'b001111111101100 : data = 16'b0000101100111110;
            15'b001111111101101 : data = 16'b0000101101000111;
            15'b001111111101110 : data = 16'b0000101101001111;
            15'b001111111101111 : data = 16'b0000101101011000;
            15'b001111111110000 : data = 16'b0000101101100000;
            15'b001111111110001 : data = 16'b0000101101101001;
            15'b001111111110010 : data = 16'b0000101101110001;
            15'b001111111110011 : data = 16'b0000101101111010;
            15'b001111111110100 : data = 16'b0000101110000010;
            15'b001111111110101 : data = 16'b0000101110001011;
            15'b001111111110110 : data = 16'b0000101110010011;
            15'b001111111110111 : data = 16'b0000101110011100;
            15'b001111111111000 : data = 16'b0000101110100100;
            15'b001111111111001 : data = 16'b0000101110101101;
            15'b001111111111010 : data = 16'b0000101110110101;
            15'b001111111111011 : data = 16'b0000101110111110;
            15'b001111111111100 : data = 16'b0000101111000111;
            15'b001111111111101 : data = 16'b0000101111001111;
            15'b001111111111110 : data = 16'b0000101111011000;
            15'b001111111111111 : data = 16'b0000101111100001;
            15'b010000000000000 : data = 16'b0000101111101001;
            15'b010000000000001 : data = 16'b0000101111110010;
            15'b010000000000010 : data = 16'b0000101111111011;
            15'b010000000000011 : data = 16'b0000110000000011;
            15'b010000000000100 : data = 16'b0000110000001100;
            15'b010000000000101 : data = 16'b0000110000010101;
            15'b010000000000110 : data = 16'b0000110000011110;
            15'b010000000000111 : data = 16'b0000110000100110;
            15'b010000000001000 : data = 16'b0000110000101111;
            15'b010000000001001 : data = 16'b0000110000111000;
            15'b010000000001010 : data = 16'b0000110001000001;
            15'b010000000001011 : data = 16'b0000110001001001;
            15'b010000000001100 : data = 16'b0000110001010010;
            15'b010000000001101 : data = 16'b0000110001011011;
            15'b010000000001110 : data = 16'b0000110001100100;
            15'b010000000001111 : data = 16'b0000110001101101;
            15'b010000000010000 : data = 16'b0000110001110110;
            15'b010000000010001 : data = 16'b0000110001111110;
            15'b010000000010010 : data = 16'b0000110010000111;
            15'b010000000010011 : data = 16'b0000110010010000;
            15'b010000000010100 : data = 16'b0000110010011001;
            15'b010000000010101 : data = 16'b0000110010100010;
            15'b010000000010110 : data = 16'b0000110010101011;
            15'b010000000010111 : data = 16'b0000110010110100;
            15'b010000000011000 : data = 16'b0000110010111101;
            15'b010000000011001 : data = 16'b0000110011000110;
            15'b010000000011010 : data = 16'b0000110011001111;
            15'b010000000011011 : data = 16'b0000110011011000;
            15'b010000000011100 : data = 16'b0000110011100001;
            15'b010000000011101 : data = 16'b0000110011101010;
            15'b010000000011110 : data = 16'b0000110011110011;
            15'b010000000011111 : data = 16'b0000110011111100;
            15'b010000000100000 : data = 16'b0000110100000101;
            15'b010000000100001 : data = 16'b0000110100001110;
            15'b010000000100010 : data = 16'b0000110100010111;
            15'b010000000100011 : data = 16'b0000110100100000;
            15'b010000000100100 : data = 16'b0000110100101001;
            15'b010000000100101 : data = 16'b0000110100110010;
            15'b010000000100110 : data = 16'b0000110100111011;
            15'b010000000100111 : data = 16'b0000110101000100;
            15'b010000000101000 : data = 16'b0000110101001110;
            15'b010000000101001 : data = 16'b0000110101010111;
            15'b010000000101010 : data = 16'b0000110101100000;
            15'b010000000101011 : data = 16'b0000110101101001;
            15'b010000000101100 : data = 16'b0000110101110010;
            15'b010000000101101 : data = 16'b0000110101111011;
            15'b010000000101110 : data = 16'b0000110110000101;
            15'b010000000101111 : data = 16'b0000110110001110;
            15'b010000000110000 : data = 16'b0000110110010111;
            15'b010000000110001 : data = 16'b0000110110100000;
            15'b010000000110010 : data = 16'b0000110110101001;
            15'b010000000110011 : data = 16'b0000110110110011;
            15'b010000000110100 : data = 16'b0000110110111100;
            15'b010000000110101 : data = 16'b0000110111000101;
            15'b010000000110110 : data = 16'b0000110111001111;
            15'b010000000110111 : data = 16'b0000110111011000;
            15'b010000000111000 : data = 16'b0000110111100001;
            15'b010000000111001 : data = 16'b0000110111101011;
            15'b010000000111010 : data = 16'b0000110111110100;
            15'b010000000111011 : data = 16'b0000110111111101;
            15'b010000000111100 : data = 16'b0000111000000111;
            15'b010000000111101 : data = 16'b0000111000010000;
            15'b010000000111110 : data = 16'b0000111000011001;
            15'b010000000111111 : data = 16'b0000111000100011;
            15'b010000001000000 : data = 16'b0000111000101100;
            15'b010000001000001 : data = 16'b0000111000110110;
            15'b010000001000010 : data = 16'b0000111000111111;
            15'b010000001000011 : data = 16'b0000111001001000;
            15'b010000001000100 : data = 16'b0000111001010010;
            15'b010000001000101 : data = 16'b0000111001011011;
            15'b010000001000110 : data = 16'b0000111001100101;
            15'b010000001000111 : data = 16'b0000111001101110;
            15'b010000001001000 : data = 16'b0000111001111000;
            15'b010000001001001 : data = 16'b0000111010000001;
            15'b010000001001010 : data = 16'b0000111010001011;
            15'b010000001001011 : data = 16'b0000111010010100;
            15'b010000001001100 : data = 16'b0000111010011110;
            15'b010000001001101 : data = 16'b0000111010101000;
            15'b010000001001110 : data = 16'b0000111010110001;
            15'b010000001001111 : data = 16'b0000111010111011;
            15'b010000001010000 : data = 16'b0000111011000100;
            15'b010000001010001 : data = 16'b0000111011001110;
            15'b010000001010010 : data = 16'b0000111011011000;
            15'b010000001010011 : data = 16'b0000111011100001;
            15'b010000001010100 : data = 16'b0000111011101011;
            15'b010000001010101 : data = 16'b0000111011110100;
            15'b010000001010110 : data = 16'b0000111011111110;
            15'b010000001010111 : data = 16'b0000111100001000;
            15'b010000001011000 : data = 16'b0000111100010001;
            15'b010000001011001 : data = 16'b0000111100011011;
            15'b010000001011010 : data = 16'b0000111100100101;
            15'b010000001011011 : data = 16'b0000111100101111;
            15'b010000001011100 : data = 16'b0000111100111000;
            15'b010000001011101 : data = 16'b0000111101000010;
            15'b010000001011110 : data = 16'b0000111101001100;
            15'b010000001011111 : data = 16'b0000111101010110;
            15'b010000001100000 : data = 16'b0000111101011111;
            15'b010000001100001 : data = 16'b0000111101101001;
            15'b010000001100010 : data = 16'b0000111101110011;
            15'b010000001100011 : data = 16'b0000111101111101;
            15'b010000001100100 : data = 16'b0000111110000111;
            15'b010000001100101 : data = 16'b0000111110010000;
            15'b010000001100110 : data = 16'b0000111110011010;
            15'b010000001100111 : data = 16'b0000111110100100;
            15'b010000001101000 : data = 16'b0000111110101110;
            15'b010000001101001 : data = 16'b0000111110111000;
            15'b010000001101010 : data = 16'b0000111111000010;
            15'b010000001101011 : data = 16'b0000111111001100;
            15'b010000001101100 : data = 16'b0000111111010110;
            15'b010000001101101 : data = 16'b0000111111011111;
            15'b010000001101110 : data = 16'b0000111111101001;
            15'b010000001101111 : data = 16'b0000111111110011;
            15'b010000001110000 : data = 16'b0000111111111101;
            15'b010000001110001 : data = 16'b0001000000000111;
            15'b010000001110010 : data = 16'b0001000000010001;
            15'b010000001110011 : data = 16'b0001000000011011;
            15'b010000001110100 : data = 16'b0001000000100101;
            15'b010000001110101 : data = 16'b0001000000101111;
            15'b010000001110110 : data = 16'b0001000000111001;
            15'b010000001110111 : data = 16'b0001000001000011;
            15'b010000001111000 : data = 16'b0001000001001101;
            15'b010000001111001 : data = 16'b0001000001010111;
            15'b010000001111010 : data = 16'b0001000001100010;
            15'b010000001111011 : data = 16'b0001000001101100;
            15'b010000001111100 : data = 16'b0001000001110110;
            15'b010000001111101 : data = 16'b0001000010000000;
            15'b010000001111110 : data = 16'b0001000010001010;
            15'b010000001111111 : data = 16'b0001000010010100;
            15'b010000010000000 : data = 16'b0001000010011110;
            15'b010000010000001 : data = 16'b0001000010101000;
            15'b010000010000010 : data = 16'b0001000010110011;
            15'b010000010000011 : data = 16'b0001000010111101;
            15'b010000010000100 : data = 16'b0001000011000111;
            15'b010000010000101 : data = 16'b0001000011010001;
            15'b010000010000110 : data = 16'b0001000011011011;
            15'b010000010000111 : data = 16'b0001000011100101;
            15'b010000010001000 : data = 16'b0001000011110000;
            15'b010000010001001 : data = 16'b0001000011111010;
            15'b010000010001010 : data = 16'b0001000100000100;
            15'b010000010001011 : data = 16'b0001000100001110;
            15'b010000010001100 : data = 16'b0001000100011001;
            15'b010000010001101 : data = 16'b0001000100100011;
            15'b010000010001110 : data = 16'b0001000100101101;
            15'b010000010001111 : data = 16'b0001000100111000;
            15'b010000010010000 : data = 16'b0001000101000010;
            15'b010000010010001 : data = 16'b0001000101001100;
            15'b010000010010010 : data = 16'b0001000101010111;
            15'b010000010010011 : data = 16'b0001000101100001;
            15'b010000010010100 : data = 16'b0001000101101011;
            15'b010000010010101 : data = 16'b0001000101110110;
            15'b010000010010110 : data = 16'b0001000110000000;
            15'b010000010010111 : data = 16'b0001000110001010;
            15'b010000010011000 : data = 16'b0001000110010101;
            15'b010000010011001 : data = 16'b0001000110011111;
            15'b010000010011010 : data = 16'b0001000110101010;
            15'b010000010011011 : data = 16'b0001000110110100;
            15'b010000010011100 : data = 16'b0001000110111111;
            15'b010000010011101 : data = 16'b0001000111001001;
            15'b010000010011110 : data = 16'b0001000111010100;
            15'b010000010011111 : data = 16'b0001000111011110;
            15'b010000010100000 : data = 16'b0001000111101001;
            15'b010000010100001 : data = 16'b0001000111110011;
            15'b010000010100010 : data = 16'b0001000111111110;
            15'b010000010100011 : data = 16'b0001001000001000;
            15'b010000010100100 : data = 16'b0001001000010011;
            15'b010000010100101 : data = 16'b0001001000011101;
            15'b010000010100110 : data = 16'b0001001000101000;
            15'b010000010100111 : data = 16'b0001001000110010;
            15'b010000010101000 : data = 16'b0001001000111101;
            15'b010000010101001 : data = 16'b0001001001001000;
            15'b010000010101010 : data = 16'b0001001001010010;
            15'b010000010101011 : data = 16'b0001001001011101;
            15'b010000010101100 : data = 16'b0001001001100111;
            15'b010000010101101 : data = 16'b0001001001110010;
            15'b010000010101110 : data = 16'b0001001001111101;
            15'b010000010101111 : data = 16'b0001001010000111;
            15'b010000010110000 : data = 16'b0001001010010010;
            15'b010000010110001 : data = 16'b0001001010011101;
            15'b010000010110010 : data = 16'b0001001010100111;
            15'b010000010110011 : data = 16'b0001001010110010;
            15'b010000010110100 : data = 16'b0001001010111101;
            15'b010000010110101 : data = 16'b0001001011001000;
            15'b010000010110110 : data = 16'b0001001011010010;
            15'b010000010110111 : data = 16'b0001001011011101;
            15'b010000010111000 : data = 16'b0001001011101000;
            15'b010000010111001 : data = 16'b0001001011110011;
            15'b010000010111010 : data = 16'b0001001011111101;
            15'b010000010111011 : data = 16'b0001001100001000;
            15'b010000010111100 : data = 16'b0001001100010011;
            15'b010000010111101 : data = 16'b0001001100011110;
            15'b010000010111110 : data = 16'b0001001100101001;
            15'b010000010111111 : data = 16'b0001001100110011;
            15'b010000011000000 : data = 16'b0001001100111110;
            15'b010000011000001 : data = 16'b0001001101001001;
            15'b010000011000010 : data = 16'b0001001101010100;
            15'b010000011000011 : data = 16'b0001001101011111;
            15'b010000011000100 : data = 16'b0001001101101010;
            15'b010000011000101 : data = 16'b0001001101110101;
            15'b010000011000110 : data = 16'b0001001110000000;
            15'b010000011000111 : data = 16'b0001001110001011;
            15'b010000011001000 : data = 16'b0001001110010110;
            15'b010000011001001 : data = 16'b0001001110100000;
            15'b010000011001010 : data = 16'b0001001110101011;
            15'b010000011001011 : data = 16'b0001001110110110;
            15'b010000011001100 : data = 16'b0001001111000001;
            15'b010000011001101 : data = 16'b0001001111001100;
            15'b010000011001110 : data = 16'b0001001111010111;
            15'b010000011001111 : data = 16'b0001001111100010;
            15'b010000011010000 : data = 16'b0001001111101101;
            15'b010000011010001 : data = 16'b0001001111111000;
            15'b010000011010010 : data = 16'b0001010000000011;
            15'b010000011010011 : data = 16'b0001010000001111;
            15'b010000011010100 : data = 16'b0001010000011010;
            15'b010000011010101 : data = 16'b0001010000100101;
            15'b010000011010110 : data = 16'b0001010000110000;
            15'b010000011010111 : data = 16'b0001010000111011;
            15'b010000011011000 : data = 16'b0001010001000110;
            15'b010000011011001 : data = 16'b0001010001010001;
            15'b010000011011010 : data = 16'b0001010001011100;
            15'b010000011011011 : data = 16'b0001010001100111;
            15'b010000011011100 : data = 16'b0001010001110011;
            15'b010000011011101 : data = 16'b0001010001111110;
            15'b010000011011110 : data = 16'b0001010010001001;
            15'b010000011011111 : data = 16'b0001010010010100;
            15'b010000011100000 : data = 16'b0001010010011111;
            15'b010000011100001 : data = 16'b0001010010101011;
            15'b010000011100010 : data = 16'b0001010010110110;
            15'b010000011100011 : data = 16'b0001010011000001;
            15'b010000011100100 : data = 16'b0001010011001100;
            15'b010000011100101 : data = 16'b0001010011010111;
            15'b010000011100110 : data = 16'b0001010011100011;
            15'b010000011100111 : data = 16'b0001010011101110;
            15'b010000011101000 : data = 16'b0001010011111001;
            15'b010000011101001 : data = 16'b0001010100000101;
            15'b010000011101010 : data = 16'b0001010100010000;
            15'b010000011101011 : data = 16'b0001010100011011;
            15'b010000011101100 : data = 16'b0001010100100111;
            15'b010000011101101 : data = 16'b0001010100110010;
            15'b010000011101110 : data = 16'b0001010100111101;
            15'b010000011101111 : data = 16'b0001010101001001;
            15'b010000011110000 : data = 16'b0001010101010100;
            15'b010000011110001 : data = 16'b0001010101011111;
            15'b010000011110010 : data = 16'b0001010101101011;
            15'b010000011110011 : data = 16'b0001010101110110;
            15'b010000011110100 : data = 16'b0001010110000010;
            15'b010000011110101 : data = 16'b0001010110001101;
            15'b010000011110110 : data = 16'b0001010110011000;
            15'b010000011110111 : data = 16'b0001010110100100;
            15'b010000011111000 : data = 16'b0001010110101111;
            15'b010000011111001 : data = 16'b0001010110111011;
            15'b010000011111010 : data = 16'b0001010111000110;
            15'b010000011111011 : data = 16'b0001010111010010;
            15'b010000011111100 : data = 16'b0001010111011101;
            15'b010000011111101 : data = 16'b0001010111101001;
            15'b010000011111110 : data = 16'b0001010111110100;
            15'b010000011111111 : data = 16'b0001011000000000;
            15'b010000100000000 : data = 16'b0001011000001011;
            15'b010000100000001 : data = 16'b0001011000010111;
            15'b010000100000010 : data = 16'b0001011000100011;
            15'b010000100000011 : data = 16'b0001011000101110;
            15'b010000100000100 : data = 16'b0001011000111010;
            15'b010000100000101 : data = 16'b0001011001000101;
            15'b010000100000110 : data = 16'b0001011001010001;
            15'b010000100000111 : data = 16'b0001011001011101;
            15'b010000100001000 : data = 16'b0001011001101000;
            15'b010000100001001 : data = 16'b0001011001110100;
            15'b010000100001010 : data = 16'b0001011001111111;
            15'b010000100001011 : data = 16'b0001011010001011;
            15'b010000100001100 : data = 16'b0001011010010111;
            15'b010000100001101 : data = 16'b0001011010100010;
            15'b010000100001110 : data = 16'b0001011010101110;
            15'b010000100001111 : data = 16'b0001011010111010;
            15'b010000100010000 : data = 16'b0001011011000110;
            15'b010000100010001 : data = 16'b0001011011010001;
            15'b010000100010010 : data = 16'b0001011011011101;
            15'b010000100010011 : data = 16'b0001011011101001;
            15'b010000100010100 : data = 16'b0001011011110101;
            15'b010000100010101 : data = 16'b0001011100000000;
            15'b010000100010110 : data = 16'b0001011100001100;
            15'b010000100010111 : data = 16'b0001011100011000;
            15'b010000100011000 : data = 16'b0001011100100100;
            15'b010000100011001 : data = 16'b0001011100110000;
            15'b010000100011010 : data = 16'b0001011100111011;
            15'b010000100011011 : data = 16'b0001011101000111;
            15'b010000100011100 : data = 16'b0001011101010011;
            15'b010000100011101 : data = 16'b0001011101011111;
            15'b010000100011110 : data = 16'b0001011101101011;
            15'b010000100011111 : data = 16'b0001011101110111;
            15'b010000100100000 : data = 16'b0001011110000011;
            15'b010000100100001 : data = 16'b0001011110001110;
            15'b010000100100010 : data = 16'b0001011110011010;
            15'b010000100100011 : data = 16'b0001011110100110;
            15'b010000100100100 : data = 16'b0001011110110010;
            15'b010000100100101 : data = 16'b0001011110111110;
            15'b010000100100110 : data = 16'b0001011111001010;
            15'b010000100100111 : data = 16'b0001011111010110;
            15'b010000100101000 : data = 16'b0001011111100010;
            15'b010000100101001 : data = 16'b0001011111101110;
            15'b010000100101010 : data = 16'b0001011111111010;
            15'b010000100101011 : data = 16'b0001100000000110;
            15'b010000100101100 : data = 16'b0001100000010010;
            15'b010000100101101 : data = 16'b0001100000011110;
            15'b010000100101110 : data = 16'b0001100000101010;
            15'b010000100101111 : data = 16'b0001100000110110;
            15'b010000100110000 : data = 16'b0001100001000010;
            15'b010000100110001 : data = 16'b0001100001001110;
            15'b010000100110010 : data = 16'b0001100001011010;
            15'b010000100110011 : data = 16'b0001100001100110;
            15'b010000100110100 : data = 16'b0001100001110010;
            15'b010000100110101 : data = 16'b0001100001111111;
            15'b010000100110110 : data = 16'b0001100010001011;
            15'b010000100110111 : data = 16'b0001100010010111;
            15'b010000100111000 : data = 16'b0001100010100011;
            15'b010000100111001 : data = 16'b0001100010101111;
            15'b010000100111010 : data = 16'b0001100010111011;
            15'b010000100111011 : data = 16'b0001100011000111;
            15'b010000100111100 : data = 16'b0001100011010100;
            15'b010000100111101 : data = 16'b0001100011100000;
            15'b010000100111110 : data = 16'b0001100011101100;
            15'b010000100111111 : data = 16'b0001100011111000;
            15'b010000101000000 : data = 16'b0001100100000100;
            15'b010000101000001 : data = 16'b0001100100010001;
            15'b010000101000010 : data = 16'b0001100100011101;
            15'b010000101000011 : data = 16'b0001100100101001;
            15'b010000101000100 : data = 16'b0001100100110101;
            15'b010000101000101 : data = 16'b0001100101000010;
            15'b010000101000110 : data = 16'b0001100101001110;
            15'b010000101000111 : data = 16'b0001100101011010;
            15'b010000101001000 : data = 16'b0001100101100111;
            15'b010000101001001 : data = 16'b0001100101110011;
            15'b010000101001010 : data = 16'b0001100101111111;
            15'b010000101001011 : data = 16'b0001100110001100;
            15'b010000101001100 : data = 16'b0001100110011000;
            15'b010000101001101 : data = 16'b0001100110100100;
            15'b010000101001110 : data = 16'b0001100110110001;
            15'b010000101001111 : data = 16'b0001100110111101;
            15'b010000101010000 : data = 16'b0001100111001001;
            15'b010000101010001 : data = 16'b0001100111010110;
            15'b010000101010010 : data = 16'b0001100111100010;
            15'b010000101010011 : data = 16'b0001100111101111;
            15'b010000101010100 : data = 16'b0001100111111011;
            15'b010000101010101 : data = 16'b0001101000000111;
            15'b010000101010110 : data = 16'b0001101000010100;
            15'b010000101010111 : data = 16'b0001101000100000;
            15'b010000101011000 : data = 16'b0001101000101101;
            15'b010000101011001 : data = 16'b0001101000111001;
            15'b010000101011010 : data = 16'b0001101001000110;
            15'b010000101011011 : data = 16'b0001101001010010;
            15'b010000101011100 : data = 16'b0001101001011111;
            15'b010000101011101 : data = 16'b0001101001101011;
            15'b010000101011110 : data = 16'b0001101001111000;
            15'b010000101011111 : data = 16'b0001101010000100;
            15'b010000101100000 : data = 16'b0001101010010001;
            15'b010000101100001 : data = 16'b0001101010011110;
            15'b010000101100010 : data = 16'b0001101010101010;
            15'b010000101100011 : data = 16'b0001101010110111;
            15'b010000101100100 : data = 16'b0001101011000011;
            15'b010000101100101 : data = 16'b0001101011010000;
            15'b010000101100110 : data = 16'b0001101011011100;
            15'b010000101100111 : data = 16'b0001101011101001;
            15'b010000101101000 : data = 16'b0001101011110110;
            15'b010000101101001 : data = 16'b0001101100000010;
            15'b010000101101010 : data = 16'b0001101100001111;
            15'b010000101101011 : data = 16'b0001101100011100;
            15'b010000101101100 : data = 16'b0001101100101000;
            15'b010000101101101 : data = 16'b0001101100110101;
            15'b010000101101110 : data = 16'b0001101101000010;
            15'b010000101101111 : data = 16'b0001101101001110;
            15'b010000101110000 : data = 16'b0001101101011011;
            15'b010000101110001 : data = 16'b0001101101101000;
            15'b010000101110010 : data = 16'b0001101101110101;
            15'b010000101110011 : data = 16'b0001101110000001;
            15'b010000101110100 : data = 16'b0001101110001110;
            15'b010000101110101 : data = 16'b0001101110011011;
            15'b010000101110110 : data = 16'b0001101110101000;
            15'b010000101110111 : data = 16'b0001101110110100;
            15'b010000101111000 : data = 16'b0001101111000001;
            15'b010000101111001 : data = 16'b0001101111001110;
            15'b010000101111010 : data = 16'b0001101111011011;
            15'b010000101111011 : data = 16'b0001101111101000;
            15'b010000101111100 : data = 16'b0001101111110101;
            15'b010000101111101 : data = 16'b0001110000000001;
            15'b010000101111110 : data = 16'b0001110000001110;
            15'b010000101111111 : data = 16'b0001110000011011;
            15'b010000110000000 : data = 16'b0001110000101000;
            15'b010000110000001 : data = 16'b0001110000110101;
            15'b010000110000010 : data = 16'b0001110001000010;
            15'b010000110000011 : data = 16'b0001110001001111;
            15'b010000110000100 : data = 16'b0001110001011100;
            15'b010000110000101 : data = 16'b0001110001101001;
            15'b010000110000110 : data = 16'b0001110001110101;
            15'b010000110000111 : data = 16'b0001110010000010;
            15'b010000110001000 : data = 16'b0001110010001111;
            15'b010000110001001 : data = 16'b0001110010011100;
            15'b010000110001010 : data = 16'b0001110010101001;
            15'b010000110001011 : data = 16'b0001110010110110;
            15'b010000110001100 : data = 16'b0001110011000011;
            15'b010000110001101 : data = 16'b0001110011010000;
            15'b010000110001110 : data = 16'b0001110011011101;
            15'b010000110001111 : data = 16'b0001110011101010;
            15'b010000110010000 : data = 16'b0001110011110111;
            15'b010000110010001 : data = 16'b0001110100000100;
            15'b010000110010010 : data = 16'b0001110100010010;
            15'b010000110010011 : data = 16'b0001110100011111;
            15'b010000110010100 : data = 16'b0001110100101100;
            15'b010000110010101 : data = 16'b0001110100111001;
            15'b010000110010110 : data = 16'b0001110101000110;
            15'b010000110010111 : data = 16'b0001110101010011;
            15'b010000110011000 : data = 16'b0001110101100000;
            15'b010000110011001 : data = 16'b0001110101101101;
            15'b010000110011010 : data = 16'b0001110101111010;
            15'b010000110011011 : data = 16'b0001110110001000;
            15'b010000110011100 : data = 16'b0001110110010101;
            15'b010000110011101 : data = 16'b0001110110100010;
            15'b010000110011110 : data = 16'b0001110110101111;
            15'b010000110011111 : data = 16'b0001110110111100;
            15'b010000110100000 : data = 16'b0001110111001001;
            15'b010000110100001 : data = 16'b0001110111010111;
            15'b010000110100010 : data = 16'b0001110111100100;
            15'b010000110100011 : data = 16'b0001110111110001;
            15'b010000110100100 : data = 16'b0001110111111110;
            15'b010000110100101 : data = 16'b0001111000001100;
            15'b010000110100110 : data = 16'b0001111000011001;
            15'b010000110100111 : data = 16'b0001111000100110;
            15'b010000110101000 : data = 16'b0001111000110011;
            15'b010000110101001 : data = 16'b0001111001000001;
            15'b010000110101010 : data = 16'b0001111001001110;
            15'b010000110101011 : data = 16'b0001111001011011;
            15'b010000110101100 : data = 16'b0001111001101001;
            15'b010000110101101 : data = 16'b0001111001110110;
            15'b010000110101110 : data = 16'b0001111010000011;
            15'b010000110101111 : data = 16'b0001111010010001;
            15'b010000110110000 : data = 16'b0001111010011110;
            15'b010000110110001 : data = 16'b0001111010101011;
            15'b010000110110010 : data = 16'b0001111010111001;
            15'b010000110110011 : data = 16'b0001111011000110;
            15'b010000110110100 : data = 16'b0001111011010011;
            15'b010000110110101 : data = 16'b0001111011100001;
            15'b010000110110110 : data = 16'b0001111011101110;
            15'b010000110110111 : data = 16'b0001111011111100;
            15'b010000110111000 : data = 16'b0001111100001001;
            15'b010000110111001 : data = 16'b0001111100010111;
            15'b010000110111010 : data = 16'b0001111100100100;
            15'b010000110111011 : data = 16'b0001111100110001;
            15'b010000110111100 : data = 16'b0001111100111111;
            15'b010000110111101 : data = 16'b0001111101001100;
            15'b010000110111110 : data = 16'b0001111101011010;
            15'b010000110111111 : data = 16'b0001111101100111;
            15'b010000111000000 : data = 16'b0001111101110101;
            15'b010000111000001 : data = 16'b0001111110000010;
            15'b010000111000010 : data = 16'b0001111110010000;
            15'b010000111000011 : data = 16'b0001111110011110;
            15'b010000111000100 : data = 16'b0001111110101011;
            15'b010000111000101 : data = 16'b0001111110111001;
            15'b010000111000110 : data = 16'b0001111111000110;
            15'b010000111000111 : data = 16'b0001111111010100;
            15'b010000111001000 : data = 16'b0001111111100001;
            15'b010000111001001 : data = 16'b0001111111101111;
            15'b010000111001010 : data = 16'b0001111111111101;
            15'b010000111001011 : data = 16'b0010000000001010;
            15'b010000111001100 : data = 16'b0010000000011000;
            15'b010000111001101 : data = 16'b0010000000100101;
            15'b010000111001110 : data = 16'b0010000000110011;
            15'b010000111001111 : data = 16'b0010000001000001;
            15'b010000111010000 : data = 16'b0010000001001110;
            15'b010000111010001 : data = 16'b0010000001011100;
            15'b010000111010010 : data = 16'b0010000001101010;
            15'b010000111010011 : data = 16'b0010000001111000;
            15'b010000111010100 : data = 16'b0010000010000101;
            15'b010000111010101 : data = 16'b0010000010010011;
            15'b010000111010110 : data = 16'b0010000010100001;
            15'b010000111010111 : data = 16'b0010000010101110;
            15'b010000111011000 : data = 16'b0010000010111100;
            15'b010000111011001 : data = 16'b0010000011001010;
            15'b010000111011010 : data = 16'b0010000011011000;
            15'b010000111011011 : data = 16'b0010000011100101;
            15'b010000111011100 : data = 16'b0010000011110011;
            15'b010000111011101 : data = 16'b0010000100000001;
            15'b010000111011110 : data = 16'b0010000100001111;
            15'b010000111011111 : data = 16'b0010000100011101;
            15'b010000111100000 : data = 16'b0010000100101010;
            15'b010000111100001 : data = 16'b0010000100111000;
            15'b010000111100010 : data = 16'b0010000101000110;
            15'b010000111100011 : data = 16'b0010000101010100;
            15'b010000111100100 : data = 16'b0010000101100010;
            15'b010000111100101 : data = 16'b0010000101110000;
            15'b010000111100110 : data = 16'b0010000101111110;
            15'b010000111100111 : data = 16'b0010000110001100;
            15'b010000111101000 : data = 16'b0010000110011001;
            15'b010000111101001 : data = 16'b0010000110100111;
            15'b010000111101010 : data = 16'b0010000110110101;
            15'b010000111101011 : data = 16'b0010000111000011;
            15'b010000111101100 : data = 16'b0010000111010001;
            15'b010000111101101 : data = 16'b0010000111011111;
            15'b010000111101110 : data = 16'b0010000111101101;
            15'b010000111101111 : data = 16'b0010000111111011;
            15'b010000111110000 : data = 16'b0010001000001001;
            15'b010000111110001 : data = 16'b0010001000010111;
            15'b010000111110010 : data = 16'b0010001000100101;
            15'b010000111110011 : data = 16'b0010001000110011;
            15'b010000111110100 : data = 16'b0010001001000001;
            15'b010000111110101 : data = 16'b0010001001001111;
            15'b010000111110110 : data = 16'b0010001001011101;
            15'b010000111110111 : data = 16'b0010001001101011;
            15'b010000111111000 : data = 16'b0010001001111001;
            15'b010000111111001 : data = 16'b0010001010000111;
            15'b010000111111010 : data = 16'b0010001010010101;
            15'b010000111111011 : data = 16'b0010001010100011;
            15'b010000111111100 : data = 16'b0010001010110001;
            15'b010000111111101 : data = 16'b0010001010111111;
            15'b010000111111110 : data = 16'b0010001011001110;
            15'b010000111111111 : data = 16'b0010001011011100;
            15'b010001000000000 : data = 16'b0010001011101010;
            15'b010001000000001 : data = 16'b0010001011111000;
            15'b010001000000010 : data = 16'b0010001100000110;
            15'b010001000000011 : data = 16'b0010001100010100;
            15'b010001000000100 : data = 16'b0010001100100010;
            15'b010001000000101 : data = 16'b0010001100110001;
            15'b010001000000110 : data = 16'b0010001100111111;
            15'b010001000000111 : data = 16'b0010001101001101;
            15'b010001000001000 : data = 16'b0010001101011011;
            15'b010001000001001 : data = 16'b0010001101101001;
            15'b010001000001010 : data = 16'b0010001101111000;
            15'b010001000001011 : data = 16'b0010001110000110;
            15'b010001000001100 : data = 16'b0010001110010100;
            15'b010001000001101 : data = 16'b0010001110100010;
            15'b010001000001110 : data = 16'b0010001110110001;
            15'b010001000001111 : data = 16'b0010001110111111;
            15'b010001000010000 : data = 16'b0010001111001101;
            15'b010001000010001 : data = 16'b0010001111011011;
            15'b010001000010010 : data = 16'b0010001111101010;
            15'b010001000010011 : data = 16'b0010001111111000;
            15'b010001000010100 : data = 16'b0010010000000110;
            15'b010001000010101 : data = 16'b0010010000010101;
            15'b010001000010110 : data = 16'b0010010000100011;
            15'b010001000010111 : data = 16'b0010010000110001;
            15'b010001000011000 : data = 16'b0010010001000000;
            15'b010001000011001 : data = 16'b0010010001001110;
            15'b010001000011010 : data = 16'b0010010001011100;
            15'b010001000011011 : data = 16'b0010010001101011;
            15'b010001000011100 : data = 16'b0010010001111001;
            15'b010001000011101 : data = 16'b0010010010001000;
            15'b010001000011110 : data = 16'b0010010010010110;
            15'b010001000011111 : data = 16'b0010010010100100;
            15'b010001000100000 : data = 16'b0010010010110011;
            15'b010001000100001 : data = 16'b0010010011000001;
            15'b010001000100010 : data = 16'b0010010011010000;
            15'b010001000100011 : data = 16'b0010010011011110;
            15'b010001000100100 : data = 16'b0010010011101101;
            15'b010001000100101 : data = 16'b0010010011111011;
            15'b010001000100110 : data = 16'b0010010100001010;
            15'b010001000100111 : data = 16'b0010010100011000;
            15'b010001000101000 : data = 16'b0010010100100111;
            15'b010001000101001 : data = 16'b0010010100110101;
            15'b010001000101010 : data = 16'b0010010101000100;
            15'b010001000101011 : data = 16'b0010010101010010;
            15'b010001000101100 : data = 16'b0010010101100001;
            15'b010001000101101 : data = 16'b0010010101101111;
            15'b010001000101110 : data = 16'b0010010101111110;
            15'b010001000101111 : data = 16'b0010010110001100;
            15'b010001000110000 : data = 16'b0010010110011011;
            15'b010001000110001 : data = 16'b0010010110101001;
            15'b010001000110010 : data = 16'b0010010110111000;
            15'b010001000110011 : data = 16'b0010010111000111;
            15'b010001000110100 : data = 16'b0010010111010101;
            15'b010001000110101 : data = 16'b0010010111100100;
            15'b010001000110110 : data = 16'b0010010111110010;
            15'b010001000110111 : data = 16'b0010011000000001;
            15'b010001000111000 : data = 16'b0010011000010000;
            15'b010001000111001 : data = 16'b0010011000011110;
            15'b010001000111010 : data = 16'b0010011000101101;
            15'b010001000111011 : data = 16'b0010011000111100;
            15'b010001000111100 : data = 16'b0010011001001010;
            15'b010001000111101 : data = 16'b0010011001011001;
            15'b010001000111110 : data = 16'b0010011001101000;
            15'b010001000111111 : data = 16'b0010011001110111;
            15'b010001001000000 : data = 16'b0010011010000101;
            15'b010001001000001 : data = 16'b0010011010010100;
            15'b010001001000010 : data = 16'b0010011010100011;
            15'b010001001000011 : data = 16'b0010011010110001;
            15'b010001001000100 : data = 16'b0010011011000000;
            15'b010001001000101 : data = 16'b0010011011001111;
            15'b010001001000110 : data = 16'b0010011011011110;
            15'b010001001000111 : data = 16'b0010011011101101;
            15'b010001001001000 : data = 16'b0010011011111011;
            15'b010001001001001 : data = 16'b0010011100001010;
            15'b010001001001010 : data = 16'b0010011100011001;
            15'b010001001001011 : data = 16'b0010011100101000;
            15'b010001001001100 : data = 16'b0010011100110111;
            15'b010001001001101 : data = 16'b0010011101000101;
            15'b010001001001110 : data = 16'b0010011101010100;
            15'b010001001001111 : data = 16'b0010011101100011;
            15'b010001001010000 : data = 16'b0010011101110010;
            15'b010001001010001 : data = 16'b0010011110000001;
            15'b010001001010010 : data = 16'b0010011110010000;
            15'b010001001010011 : data = 16'b0010011110011111;
            15'b010001001010100 : data = 16'b0010011110101101;
            15'b010001001010101 : data = 16'b0010011110111100;
            15'b010001001010110 : data = 16'b0010011111001011;
            15'b010001001010111 : data = 16'b0010011111011010;
            15'b010001001011000 : data = 16'b0010011111101001;
            15'b010001001011001 : data = 16'b0010011111111000;
            15'b010001001011010 : data = 16'b0010100000000111;
            15'b010001001011011 : data = 16'b0010100000010110;
            15'b010001001011100 : data = 16'b0010100000100101;
            15'b010001001011101 : data = 16'b0010100000110100;
            15'b010001001011110 : data = 16'b0010100001000011;
            15'b010001001011111 : data = 16'b0010100001010010;
            15'b010001001100000 : data = 16'b0010100001100001;
            15'b010001001100001 : data = 16'b0010100001110000;
            15'b010001001100010 : data = 16'b0010100001111111;
            15'b010001001100011 : data = 16'b0010100010001110;
            15'b010001001100100 : data = 16'b0010100010011101;
            15'b010001001100101 : data = 16'b0010100010101100;
            15'b010001001100110 : data = 16'b0010100010111011;
            15'b010001001100111 : data = 16'b0010100011001010;
            15'b010001001101000 : data = 16'b0010100011011001;
            15'b010001001101001 : data = 16'b0010100011101000;
            15'b010001001101010 : data = 16'b0010100011110111;
            15'b010001001101011 : data = 16'b0010100100000111;
            15'b010001001101100 : data = 16'b0010100100010110;
            15'b010001001101101 : data = 16'b0010100100100101;
            15'b010001001101110 : data = 16'b0010100100110100;
            15'b010001001101111 : data = 16'b0010100101000011;
            15'b010001001110000 : data = 16'b0010100101010010;
            15'b010001001110001 : data = 16'b0010100101100001;
            15'b010001001110010 : data = 16'b0010100101110001;
            15'b010001001110011 : data = 16'b0010100110000000;
            15'b010001001110100 : data = 16'b0010100110001111;
            15'b010001001110101 : data = 16'b0010100110011110;
            15'b010001001110110 : data = 16'b0010100110101101;
            15'b010001001110111 : data = 16'b0010100110111100;
            15'b010001001111000 : data = 16'b0010100111001100;
            15'b010001001111001 : data = 16'b0010100111011011;
            15'b010001001111010 : data = 16'b0010100111101010;
            15'b010001001111011 : data = 16'b0010100111111001;
            15'b010001001111100 : data = 16'b0010101000001001;
            15'b010001001111101 : data = 16'b0010101000011000;
            15'b010001001111110 : data = 16'b0010101000100111;
            15'b010001001111111 : data = 16'b0010101000110110;
            15'b010001010000000 : data = 16'b0010101001000110;
            15'b010001010000001 : data = 16'b0010101001010101;
            15'b010001010000010 : data = 16'b0010101001100100;
            15'b010001010000011 : data = 16'b0010101001110100;
            15'b010001010000100 : data = 16'b0010101010000011;
            15'b010001010000101 : data = 16'b0010101010010010;
            15'b010001010000110 : data = 16'b0010101010100010;
            15'b010001010000111 : data = 16'b0010101010110001;
            15'b010001010001000 : data = 16'b0010101011000000;
            15'b010001010001001 : data = 16'b0010101011010000;
            15'b010001010001010 : data = 16'b0010101011011111;
            15'b010001010001011 : data = 16'b0010101011101110;
            15'b010001010001100 : data = 16'b0010101011111110;
            15'b010001010001101 : data = 16'b0010101100001101;
            15'b010001010001110 : data = 16'b0010101100011101;
            15'b010001010001111 : data = 16'b0010101100101100;
            15'b010001010010000 : data = 16'b0010101100111011;
            15'b010001010010001 : data = 16'b0010101101001011;
            15'b010001010010010 : data = 16'b0010101101011010;
            15'b010001010010011 : data = 16'b0010101101101010;
            15'b010001010010100 : data = 16'b0010101101111001;
            15'b010001010010101 : data = 16'b0010101110001001;
            15'b010001010010110 : data = 16'b0010101110011000;
            15'b010001010010111 : data = 16'b0010101110101000;
            15'b010001010011000 : data = 16'b0010101110110111;
            15'b010001010011001 : data = 16'b0010101111000111;
            15'b010001010011010 : data = 16'b0010101111010110;
            15'b010001010011011 : data = 16'b0010101111100110;
            15'b010001010011100 : data = 16'b0010101111110101;
            15'b010001010011101 : data = 16'b0010110000000101;
            15'b010001010011110 : data = 16'b0010110000010100;
            15'b010001010011111 : data = 16'b0010110000100100;
            15'b010001010100000 : data = 16'b0010110000110011;
            15'b010001010100001 : data = 16'b0010110001000011;
            15'b010001010100010 : data = 16'b0010110001010010;
            15'b010001010100011 : data = 16'b0010110001100010;
            15'b010001010100100 : data = 16'b0010110001110010;
            15'b010001010100101 : data = 16'b0010110010000001;
            15'b010001010100110 : data = 16'b0010110010010001;
            15'b010001010100111 : data = 16'b0010110010100000;
            15'b010001010101000 : data = 16'b0010110010110000;
            15'b010001010101001 : data = 16'b0010110011000000;
            15'b010001010101010 : data = 16'b0010110011001111;
            15'b010001010101011 : data = 16'b0010110011011111;
            15'b010001010101100 : data = 16'b0010110011101111;
            15'b010001010101101 : data = 16'b0010110011111110;
            15'b010001010101110 : data = 16'b0010110100001110;
            15'b010001010101111 : data = 16'b0010110100011110;
            15'b010001010110000 : data = 16'b0010110100101101;
            15'b010001010110001 : data = 16'b0010110100111101;
            15'b010001010110010 : data = 16'b0010110101001101;
            15'b010001010110011 : data = 16'b0010110101011101;
            15'b010001010110100 : data = 16'b0010110101101100;
            15'b010001010110101 : data = 16'b0010110101111100;
            15'b010001010110110 : data = 16'b0010110110001100;
            15'b010001010110111 : data = 16'b0010110110011100;
            15'b010001010111000 : data = 16'b0010110110101011;
            15'b010001010111001 : data = 16'b0010110110111011;
            15'b010001010111010 : data = 16'b0010110111001011;
            15'b010001010111011 : data = 16'b0010110111011011;
            15'b010001010111100 : data = 16'b0010110111101010;
            15'b010001010111101 : data = 16'b0010110111111010;
            15'b010001010111110 : data = 16'b0010111000001010;
            15'b010001010111111 : data = 16'b0010111000011010;
            15'b010001011000000 : data = 16'b0010111000101010;
            15'b010001011000001 : data = 16'b0010111000111001;
            15'b010001011000010 : data = 16'b0010111001001001;
            15'b010001011000011 : data = 16'b0010111001011001;
            15'b010001011000100 : data = 16'b0010111001101001;
            15'b010001011000101 : data = 16'b0010111001111001;
            15'b010001011000110 : data = 16'b0010111010001001;
            15'b010001011000111 : data = 16'b0010111010011001;
            15'b010001011001000 : data = 16'b0010111010101001;
            15'b010001011001001 : data = 16'b0010111010111000;
            15'b010001011001010 : data = 16'b0010111011001000;
            15'b010001011001011 : data = 16'b0010111011011000;
            15'b010001011001100 : data = 16'b0010111011101000;
            15'b010001011001101 : data = 16'b0010111011111000;
            15'b010001011001110 : data = 16'b0010111100001000;
            15'b010001011001111 : data = 16'b0010111100011000;
            15'b010001011010000 : data = 16'b0010111100101000;
            15'b010001011010001 : data = 16'b0010111100111000;
            15'b010001011010010 : data = 16'b0010111101001000;
            15'b010001011010011 : data = 16'b0010111101011000;
            15'b010001011010100 : data = 16'b0010111101101000;
            15'b010001011010101 : data = 16'b0010111101111000;
            15'b010001011010110 : data = 16'b0010111110001000;
            15'b010001011010111 : data = 16'b0010111110011000;
            15'b010001011011000 : data = 16'b0010111110101000;
            15'b010001011011001 : data = 16'b0010111110111000;
            15'b010001011011010 : data = 16'b0010111111001000;
            15'b010001011011011 : data = 16'b0010111111011000;
            15'b010001011011100 : data = 16'b0010111111101000;
            15'b010001011011101 : data = 16'b0010111111111000;
            15'b010001011011110 : data = 16'b0011000000001000;
            15'b010001011011111 : data = 16'b0011000000011000;
            15'b010001011100000 : data = 16'b0011000000101000;
            15'b010001011100001 : data = 16'b0011000000111001;
            15'b010001011100010 : data = 16'b0011000001001001;
            15'b010001011100011 : data = 16'b0011000001011001;
            15'b010001011100100 : data = 16'b0011000001101001;
            15'b010001011100101 : data = 16'b0011000001111001;
            15'b010001011100110 : data = 16'b0011000010001001;
            15'b010001011100111 : data = 16'b0011000010011001;
            15'b010001011101000 : data = 16'b0011000010101001;
            15'b010001011101001 : data = 16'b0011000010111010;
            15'b010001011101010 : data = 16'b0011000011001010;
            15'b010001011101011 : data = 16'b0011000011011010;
            15'b010001011101100 : data = 16'b0011000011101010;
            15'b010001011101101 : data = 16'b0011000011111010;
            15'b010001011101110 : data = 16'b0011000100001010;
            15'b010001011101111 : data = 16'b0011000100011011;
            15'b010001011110000 : data = 16'b0011000100101011;
            15'b010001011110001 : data = 16'b0011000100111011;
            15'b010001011110010 : data = 16'b0011000101001011;
            15'b010001011110011 : data = 16'b0011000101011100;
            15'b010001011110100 : data = 16'b0011000101101100;
            15'b010001011110101 : data = 16'b0011000101111100;
            15'b010001011110110 : data = 16'b0011000110001100;
            15'b010001011110111 : data = 16'b0011000110011101;
            15'b010001011111000 : data = 16'b0011000110101101;
            15'b010001011111001 : data = 16'b0011000110111101;
            15'b010001011111010 : data = 16'b0011000111001110;
            15'b010001011111011 : data = 16'b0011000111011110;
            15'b010001011111100 : data = 16'b0011000111101110;
            15'b010001011111101 : data = 16'b0011000111111110;
            15'b010001011111110 : data = 16'b0011001000001111;
            15'b010001011111111 : data = 16'b0011001000011111;
            15'b010001100000000 : data = 16'b0011001000101111;
            15'b010001100000001 : data = 16'b0011001001000000;
            15'b010001100000010 : data = 16'b0011001001010000;
            15'b010001100000011 : data = 16'b0011001001100001;
            15'b010001100000100 : data = 16'b0011001001110001;
            15'b010001100000101 : data = 16'b0011001010000001;
            15'b010001100000110 : data = 16'b0011001010010010;
            15'b010001100000111 : data = 16'b0011001010100010;
            15'b010001100001000 : data = 16'b0011001010110010;
            15'b010001100001001 : data = 16'b0011001011000011;
            15'b010001100001010 : data = 16'b0011001011010011;
            15'b010001100001011 : data = 16'b0011001011100100;
            15'b010001100001100 : data = 16'b0011001011110100;
            15'b010001100001101 : data = 16'b0011001100000101;
            15'b010001100001110 : data = 16'b0011001100010101;
            15'b010001100001111 : data = 16'b0011001100100110;
            15'b010001100010000 : data = 16'b0011001100110110;
            15'b010001100010001 : data = 16'b0011001101000110;
            15'b010001100010010 : data = 16'b0011001101010111;
            15'b010001100010011 : data = 16'b0011001101100111;
            15'b010001100010100 : data = 16'b0011001101111000;
            15'b010001100010101 : data = 16'b0011001110001000;
            15'b010001100010110 : data = 16'b0011001110011001;
            15'b010001100010111 : data = 16'b0011001110101001;
            15'b010001100011000 : data = 16'b0011001110111010;
            15'b010001100011001 : data = 16'b0011001111001011;
            15'b010001100011010 : data = 16'b0011001111011011;
            15'b010001100011011 : data = 16'b0011001111101100;
            15'b010001100011100 : data = 16'b0011001111111100;
            15'b010001100011101 : data = 16'b0011010000001101;
            15'b010001100011110 : data = 16'b0011010000011101;
            15'b010001100011111 : data = 16'b0011010000101110;
            15'b010001100100000 : data = 16'b0011010000111111;
            15'b010001100100001 : data = 16'b0011010001001111;
            15'b010001100100010 : data = 16'b0011010001100000;
            15'b010001100100011 : data = 16'b0011010001110000;
            15'b010001100100100 : data = 16'b0011010010000001;
            15'b010001100100101 : data = 16'b0011010010010010;
            15'b010001100100110 : data = 16'b0011010010100010;
            15'b010001100100111 : data = 16'b0011010010110011;
            15'b010001100101000 : data = 16'b0011010011000100;
            15'b010001100101001 : data = 16'b0011010011010100;
            15'b010001100101010 : data = 16'b0011010011100101;
            15'b010001100101011 : data = 16'b0011010011110110;
            15'b010001100101100 : data = 16'b0011010100000110;
            15'b010001100101101 : data = 16'b0011010100010111;
            15'b010001100101110 : data = 16'b0011010100101000;
            15'b010001100101111 : data = 16'b0011010100111000;
            15'b010001100110000 : data = 16'b0011010101001001;
            15'b010001100110001 : data = 16'b0011010101011010;
            15'b010001100110010 : data = 16'b0011010101101010;
            15'b010001100110011 : data = 16'b0011010101111011;
            15'b010001100110100 : data = 16'b0011010110001100;
            15'b010001100110101 : data = 16'b0011010110011101;
            15'b010001100110110 : data = 16'b0011010110101101;
            15'b010001100110111 : data = 16'b0011010110111110;
            15'b010001100111000 : data = 16'b0011010111001111;
            15'b010001100111001 : data = 16'b0011010111100000;
            15'b010001100111010 : data = 16'b0011010111110001;
            15'b010001100111011 : data = 16'b0011011000000001;
            15'b010001100111100 : data = 16'b0011011000010010;
            15'b010001100111101 : data = 16'b0011011000100011;
            15'b010001100111110 : data = 16'b0011011000110100;
            15'b010001100111111 : data = 16'b0011011001000101;
            15'b010001101000000 : data = 16'b0011011001010101;
            15'b010001101000001 : data = 16'b0011011001100110;
            15'b010001101000010 : data = 16'b0011011001110111;
            15'b010001101000011 : data = 16'b0011011010001000;
            15'b010001101000100 : data = 16'b0011011010011001;
            15'b010001101000101 : data = 16'b0011011010101010;
            15'b010001101000110 : data = 16'b0011011010111011;
            15'b010001101000111 : data = 16'b0011011011001100;
            15'b010001101001000 : data = 16'b0011011011011100;
            15'b010001101001001 : data = 16'b0011011011101101;
            15'b010001101001010 : data = 16'b0011011011111110;
            15'b010001101001011 : data = 16'b0011011100001111;
            15'b010001101001100 : data = 16'b0011011100100000;
            15'b010001101001101 : data = 16'b0011011100110001;
            15'b010001101001110 : data = 16'b0011011101000010;
            15'b010001101001111 : data = 16'b0011011101010011;
            15'b010001101010000 : data = 16'b0011011101100100;
            15'b010001101010001 : data = 16'b0011011101110101;
            15'b010001101010010 : data = 16'b0011011110000110;
            15'b010001101010011 : data = 16'b0011011110010111;
            15'b010001101010100 : data = 16'b0011011110101000;
            15'b010001101010101 : data = 16'b0011011110111001;
            15'b010001101010110 : data = 16'b0011011111001010;
            15'b010001101010111 : data = 16'b0011011111011011;
            15'b010001101011000 : data = 16'b0011011111101100;
            15'b010001101011001 : data = 16'b0011011111111101;
            15'b010001101011010 : data = 16'b0011100000001110;
            15'b010001101011011 : data = 16'b0011100000011111;
            15'b010001101011100 : data = 16'b0011100000110000;
            15'b010001101011101 : data = 16'b0011100001000001;
            15'b010001101011110 : data = 16'b0011100001010010;
            15'b010001101011111 : data = 16'b0011100001100011;
            15'b010001101100000 : data = 16'b0011100001110100;
            15'b010001101100001 : data = 16'b0011100010000101;
            15'b010001101100010 : data = 16'b0011100010010110;
            15'b010001101100011 : data = 16'b0011100010100111;
            15'b010001101100100 : data = 16'b0011100010111000;
            15'b010001101100101 : data = 16'b0011100011001001;
            15'b010001101100110 : data = 16'b0011100011011011;
            15'b010001101100111 : data = 16'b0011100011101100;
            15'b010001101101000 : data = 16'b0011100011111101;
            15'b010001101101001 : data = 16'b0011100100001110;
            15'b010001101101010 : data = 16'b0011100100011111;
            15'b010001101101011 : data = 16'b0011100100110000;
            15'b010001101101100 : data = 16'b0011100101000001;
            15'b010001101101101 : data = 16'b0011100101010011;
            15'b010001101101110 : data = 16'b0011100101100100;
            15'b010001101101111 : data = 16'b0011100101110101;
            15'b010001101110000 : data = 16'b0011100110000110;
            15'b010001101110001 : data = 16'b0011100110010111;
            15'b010001101110010 : data = 16'b0011100110101000;
            15'b010001101110011 : data = 16'b0011100110111010;
            15'b010001101110100 : data = 16'b0011100111001011;
            15'b010001101110101 : data = 16'b0011100111011100;
            15'b010001101110110 : data = 16'b0011100111101101;
            15'b010001101110111 : data = 16'b0011100111111111;
            15'b010001101111000 : data = 16'b0011101000010000;
            15'b010001101111001 : data = 16'b0011101000100001;
            15'b010001101111010 : data = 16'b0011101000110010;
            15'b010001101111011 : data = 16'b0011101001000100;
            15'b010001101111100 : data = 16'b0011101001010101;
            15'b010001101111101 : data = 16'b0011101001100110;
            15'b010001101111110 : data = 16'b0011101001110111;
            15'b010001101111111 : data = 16'b0011101010001001;
            15'b010001110000000 : data = 16'b0011101010011010;
            15'b010001110000001 : data = 16'b0011101010101011;
            15'b010001110000010 : data = 16'b0011101010111101;
            15'b010001110000011 : data = 16'b0011101011001110;
            15'b010001110000100 : data = 16'b0011101011011111;
            15'b010001110000101 : data = 16'b0011101011110001;
            15'b010001110000110 : data = 16'b0011101100000010;
            15'b010001110000111 : data = 16'b0011101100010011;
            15'b010001110001000 : data = 16'b0011101100100101;
            15'b010001110001001 : data = 16'b0011101100110110;
            15'b010001110001010 : data = 16'b0011101101000111;
            15'b010001110001011 : data = 16'b0011101101011001;
            15'b010001110001100 : data = 16'b0011101101101010;
            15'b010001110001101 : data = 16'b0011101101111011;
            15'b010001110001110 : data = 16'b0011101110001101;
            15'b010001110001111 : data = 16'b0011101110011110;
            15'b010001110010000 : data = 16'b0011101110110000;
            15'b010001110010001 : data = 16'b0011101111000001;
            15'b010001110010010 : data = 16'b0011101111010010;
            15'b010001110010011 : data = 16'b0011101111100100;
            15'b010001110010100 : data = 16'b0011101111110101;
            15'b010001110010101 : data = 16'b0011110000000111;
            15'b010001110010110 : data = 16'b0011110000011000;
            15'b010001110010111 : data = 16'b0011110000101010;
            15'b010001110011000 : data = 16'b0011110000111011;
            15'b010001110011001 : data = 16'b0011110001001101;
            15'b010001110011010 : data = 16'b0011110001011110;
            15'b010001110011011 : data = 16'b0011110001110000;
            15'b010001110011100 : data = 16'b0011110010000001;
            15'b010001110011101 : data = 16'b0011110010010011;
            15'b010001110011110 : data = 16'b0011110010100100;
            15'b010001110011111 : data = 16'b0011110010110110;
            15'b010001110100000 : data = 16'b0011110011000111;
            15'b010001110100001 : data = 16'b0011110011011001;
            15'b010001110100010 : data = 16'b0011110011101010;
            15'b010001110100011 : data = 16'b0011110011111100;
            15'b010001110100100 : data = 16'b0011110100001101;
            15'b010001110100101 : data = 16'b0011110100011111;
            15'b010001110100110 : data = 16'b0011110100110000;
            15'b010001110100111 : data = 16'b0011110101000010;
            15'b010001110101000 : data = 16'b0011110101010011;
            15'b010001110101001 : data = 16'b0011110101100101;
            15'b010001110101010 : data = 16'b0011110101110111;
            15'b010001110101011 : data = 16'b0011110110001000;
            15'b010001110101100 : data = 16'b0011110110011010;
            15'b010001110101101 : data = 16'b0011110110101011;
            15'b010001110101110 : data = 16'b0011110110111101;
            15'b010001110101111 : data = 16'b0011110111001111;
            15'b010001110110000 : data = 16'b0011110111100000;
            15'b010001110110001 : data = 16'b0011110111110010;
            15'b010001110110010 : data = 16'b0011111000000100;
            15'b010001110110011 : data = 16'b0011111000010101;
            15'b010001110110100 : data = 16'b0011111000100111;
            15'b010001110110101 : data = 16'b0011111000111001;
            15'b010001110110110 : data = 16'b0011111001001010;
            15'b010001110110111 : data = 16'b0011111001011100;
            15'b010001110111000 : data = 16'b0011111001101110;
            15'b010001110111001 : data = 16'b0011111001111111;
            15'b010001110111010 : data = 16'b0011111010010001;
            15'b010001110111011 : data = 16'b0011111010100011;
            15'b010001110111100 : data = 16'b0011111010110100;
            15'b010001110111101 : data = 16'b0011111011000110;
            15'b010001110111110 : data = 16'b0011111011011000;
            15'b010001110111111 : data = 16'b0011111011101001;
            15'b010001111000000 : data = 16'b0011111011111011;
            15'b010001111000001 : data = 16'b0011111100001101;
            15'b010001111000010 : data = 16'b0011111100011111;
            15'b010001111000011 : data = 16'b0011111100110000;
            15'b010001111000100 : data = 16'b0011111101000010;
            15'b010001111000101 : data = 16'b0011111101010100;
            15'b010001111000110 : data = 16'b0011111101100110;
            15'b010001111000111 : data = 16'b0011111101110111;
            15'b010001111001000 : data = 16'b0011111110001001;
            15'b010001111001001 : data = 16'b0011111110011011;
            15'b010001111001010 : data = 16'b0011111110101101;
            15'b010001111001011 : data = 16'b0011111110111111;
            15'b010001111001100 : data = 16'b0011111111010000;
            15'b010001111001101 : data = 16'b0011111111100010;
            15'b010001111001110 : data = 16'b0011111111110100;
            15'b010001111001111 : data = 16'b0100000000000110;
            15'b010001111010000 : data = 16'b0100000000011000;
            15'b010001111010001 : data = 16'b0100000000101010;
            15'b010001111010010 : data = 16'b0100000000111011;
            15'b010001111010011 : data = 16'b0100000001001101;
            15'b010001111010100 : data = 16'b0100000001011111;
            15'b010001111010101 : data = 16'b0100000001110001;
            15'b010001111010110 : data = 16'b0100000010000011;
            15'b010001111010111 : data = 16'b0100000010010101;
            15'b010001111011000 : data = 16'b0100000010100111;
            15'b010001111011001 : data = 16'b0100000010111001;
            15'b010001111011010 : data = 16'b0100000011001010;
            15'b010001111011011 : data = 16'b0100000011011100;
            15'b010001111011100 : data = 16'b0100000011101110;
            15'b010001111011101 : data = 16'b0100000100000000;
            15'b010001111011110 : data = 16'b0100000100010010;
            15'b010001111011111 : data = 16'b0100000100100100;
            15'b010001111100000 : data = 16'b0100000100110110;
            15'b010001111100001 : data = 16'b0100000101001000;
            15'b010001111100010 : data = 16'b0100000101011010;
            15'b010001111100011 : data = 16'b0100000101101100;
            15'b010001111100100 : data = 16'b0100000101111110;
            15'b010001111100101 : data = 16'b0100000110010000;
            15'b010001111100110 : data = 16'b0100000110100010;
            15'b010001111100111 : data = 16'b0100000110110100;
            15'b010001111101000 : data = 16'b0100000111000110;
            15'b010001111101001 : data = 16'b0100000111011000;
            15'b010001111101010 : data = 16'b0100000111101010;
            15'b010001111101011 : data = 16'b0100000111111100;
            15'b010001111101100 : data = 16'b0100001000001110;
            15'b010001111101101 : data = 16'b0100001000100000;
            15'b010001111101110 : data = 16'b0100001000110010;
            15'b010001111101111 : data = 16'b0100001001000100;
            15'b010001111110000 : data = 16'b0100001001010110;
            15'b010001111110001 : data = 16'b0100001001101000;
            15'b010001111110010 : data = 16'b0100001001111010;
            15'b010001111110011 : data = 16'b0100001010001100;
            15'b010001111110100 : data = 16'b0100001010011110;
            15'b010001111110101 : data = 16'b0100001010110000;
            15'b010001111110110 : data = 16'b0100001011000010;
            15'b010001111110111 : data = 16'b0100001011010100;
            15'b010001111111000 : data = 16'b0100001011100110;
            15'b010001111111001 : data = 16'b0100001011111001;
            15'b010001111111010 : data = 16'b0100001100001011;
            15'b010001111111011 : data = 16'b0100001100011101;
            15'b010001111111100 : data = 16'b0100001100101111;
            15'b010001111111101 : data = 16'b0100001101000001;
            15'b010001111111110 : data = 16'b0100001101010011;
            15'b010001111111111 : data = 16'b0100001101100101;
            15'b010010000000000 : data = 16'b0100001101110111;
            15'b010010000000001 : data = 16'b0100001110001001;
            15'b010010000000010 : data = 16'b0100001110011100;
            15'b010010000000011 : data = 16'b0100001110101110;
            15'b010010000000100 : data = 16'b0100001111000000;
            15'b010010000000101 : data = 16'b0100001111010010;
            15'b010010000000110 : data = 16'b0100001111100100;
            15'b010010000000111 : data = 16'b0100001111110110;
            15'b010010000001000 : data = 16'b0100010000001001;
            15'b010010000001001 : data = 16'b0100010000011011;
            15'b010010000001010 : data = 16'b0100010000101101;
            15'b010010000001011 : data = 16'b0100010000111111;
            15'b010010000001100 : data = 16'b0100010001010001;
            15'b010010000001101 : data = 16'b0100010001100100;
            15'b010010000001110 : data = 16'b0100010001110110;
            15'b010010000001111 : data = 16'b0100010010001000;
            15'b010010000010000 : data = 16'b0100010010011010;
            15'b010010000010001 : data = 16'b0100010010101101;
            15'b010010000010010 : data = 16'b0100010010111111;
            15'b010010000010011 : data = 16'b0100010011010001;
            15'b010010000010100 : data = 16'b0100010011100011;
            15'b010010000010101 : data = 16'b0100010011110110;
            15'b010010000010110 : data = 16'b0100010100001000;
            15'b010010000010111 : data = 16'b0100010100011010;
            15'b010010000011000 : data = 16'b0100010100101100;
            15'b010010000011001 : data = 16'b0100010100111111;
            15'b010010000011010 : data = 16'b0100010101010001;
            15'b010010000011011 : data = 16'b0100010101100011;
            15'b010010000011100 : data = 16'b0100010101110110;
            15'b010010000011101 : data = 16'b0100010110001000;
            15'b010010000011110 : data = 16'b0100010110011010;
            15'b010010000011111 : data = 16'b0100010110101101;
            15'b010010000100000 : data = 16'b0100010110111111;
            15'b010010000100001 : data = 16'b0100010111010001;
            15'b010010000100010 : data = 16'b0100010111100100;
            15'b010010000100011 : data = 16'b0100010111110110;
            15'b010010000100100 : data = 16'b0100011000001000;
            15'b010010000100101 : data = 16'b0100011000011011;
            15'b010010000100110 : data = 16'b0100011000101101;
            15'b010010000100111 : data = 16'b0100011000111111;
            15'b010010000101000 : data = 16'b0100011001010010;
            15'b010010000101001 : data = 16'b0100011001100100;
            15'b010010000101010 : data = 16'b0100011001110111;
            15'b010010000101011 : data = 16'b0100011010001001;
            15'b010010000101100 : data = 16'b0100011010011011;
            15'b010010000101101 : data = 16'b0100011010101110;
            15'b010010000101110 : data = 16'b0100011011000000;
            15'b010010000101111 : data = 16'b0100011011010011;
            15'b010010000110000 : data = 16'b0100011011100101;
            15'b010010000110001 : data = 16'b0100011011110111;
            15'b010010000110010 : data = 16'b0100011100001010;
            15'b010010000110011 : data = 16'b0100011100011100;
            15'b010010000110100 : data = 16'b0100011100101111;
            15'b010010000110101 : data = 16'b0100011101000001;
            15'b010010000110110 : data = 16'b0100011101010100;
            15'b010010000110111 : data = 16'b0100011101100110;
            15'b010010000111000 : data = 16'b0100011101111001;
            15'b010010000111001 : data = 16'b0100011110001011;
            15'b010010000111010 : data = 16'b0100011110011110;
            15'b010010000111011 : data = 16'b0100011110110000;
            15'b010010000111100 : data = 16'b0100011111000011;
            15'b010010000111101 : data = 16'b0100011111010101;
            15'b010010000111110 : data = 16'b0100011111101000;
            15'b010010000111111 : data = 16'b0100011111111010;
            15'b010010001000000 : data = 16'b0100100000001101;
            15'b010010001000001 : data = 16'b0100100000011111;
            15'b010010001000010 : data = 16'b0100100000110010;
            15'b010010001000011 : data = 16'b0100100001000100;
            15'b010010001000100 : data = 16'b0100100001010111;
            15'b010010001000101 : data = 16'b0100100001101001;
            15'b010010001000110 : data = 16'b0100100001111100;
            15'b010010001000111 : data = 16'b0100100010001110;
            15'b010010001001000 : data = 16'b0100100010100001;
            15'b010010001001001 : data = 16'b0100100010110011;
            15'b010010001001010 : data = 16'b0100100011000110;
            15'b010010001001011 : data = 16'b0100100011011001;
            15'b010010001001100 : data = 16'b0100100011101011;
            15'b010010001001101 : data = 16'b0100100011111110;
            15'b010010001001110 : data = 16'b0100100100010000;
            15'b010010001001111 : data = 16'b0100100100100011;
            15'b010010001010000 : data = 16'b0100100100110110;
            15'b010010001010001 : data = 16'b0100100101001000;
            15'b010010001010010 : data = 16'b0100100101011011;
            15'b010010001010011 : data = 16'b0100100101101101;
            15'b010010001010100 : data = 16'b0100100110000000;
            15'b010010001010101 : data = 16'b0100100110010011;
            15'b010010001010110 : data = 16'b0100100110100101;
            15'b010010001010111 : data = 16'b0100100110111000;
            15'b010010001011000 : data = 16'b0100100111001011;
            15'b010010001011001 : data = 16'b0100100111011101;
            15'b010010001011010 : data = 16'b0100100111110000;
            15'b010010001011011 : data = 16'b0100101000000011;
            15'b010010001011100 : data = 16'b0100101000010101;
            15'b010010001011101 : data = 16'b0100101000101000;
            15'b010010001011110 : data = 16'b0100101000111011;
            15'b010010001011111 : data = 16'b0100101001001101;
            15'b010010001100000 : data = 16'b0100101001100000;
            15'b010010001100001 : data = 16'b0100101001110011;
            15'b010010001100010 : data = 16'b0100101010000101;
            15'b010010001100011 : data = 16'b0100101010011000;
            15'b010010001100100 : data = 16'b0100101010101011;
            15'b010010001100101 : data = 16'b0100101010111101;
            15'b010010001100110 : data = 16'b0100101011010000;
            15'b010010001100111 : data = 16'b0100101011100011;
            15'b010010001101000 : data = 16'b0100101011110110;
            15'b010010001101001 : data = 16'b0100101100001000;
            15'b010010001101010 : data = 16'b0100101100011011;
            15'b010010001101011 : data = 16'b0100101100101110;
            15'b010010001101100 : data = 16'b0100101101000001;
            15'b010010001101101 : data = 16'b0100101101010011;
            15'b010010001101110 : data = 16'b0100101101100110;
            15'b010010001101111 : data = 16'b0100101101111001;
            15'b010010001110000 : data = 16'b0100101110001100;
            15'b010010001110001 : data = 16'b0100101110011111;
            15'b010010001110010 : data = 16'b0100101110110001;
            15'b010010001110011 : data = 16'b0100101111000100;
            15'b010010001110100 : data = 16'b0100101111010111;
            15'b010010001110101 : data = 16'b0100101111101010;
            15'b010010001110110 : data = 16'b0100101111111101;
            15'b010010001110111 : data = 16'b0100110000001111;
            15'b010010001111000 : data = 16'b0100110000100010;
            15'b010010001111001 : data = 16'b0100110000110101;
            15'b010010001111010 : data = 16'b0100110001001000;
            15'b010010001111011 : data = 16'b0100110001011011;
            15'b010010001111100 : data = 16'b0100110001101101;
            15'b010010001111101 : data = 16'b0100110010000000;
            15'b010010001111110 : data = 16'b0100110010010011;
            15'b010010001111111 : data = 16'b0100110010100110;
            15'b010010010000000 : data = 16'b0100110010111001;
            15'b010010010000001 : data = 16'b0100110011001100;
            15'b010010010000010 : data = 16'b0100110011011111;
            15'b010010010000011 : data = 16'b0100110011110001;
            15'b010010010000100 : data = 16'b0100110100000100;
            15'b010010010000101 : data = 16'b0100110100010111;
            15'b010010010000110 : data = 16'b0100110100101010;
            15'b010010010000111 : data = 16'b0100110100111101;
            15'b010010010001000 : data = 16'b0100110101010000;
            15'b010010010001001 : data = 16'b0100110101100011;
            15'b010010010001010 : data = 16'b0100110101110110;
            15'b010010010001011 : data = 16'b0100110110001001;
            15'b010010010001100 : data = 16'b0100110110011100;
            15'b010010010001101 : data = 16'b0100110110101111;
            15'b010010010001110 : data = 16'b0100110111000001;
            15'b010010010001111 : data = 16'b0100110111010100;
            15'b010010010010000 : data = 16'b0100110111100111;
            15'b010010010010001 : data = 16'b0100110111111010;
            15'b010010010010010 : data = 16'b0100111000001101;
            15'b010010010010011 : data = 16'b0100111000100000;
            15'b010010010010100 : data = 16'b0100111000110011;
            15'b010010010010101 : data = 16'b0100111001000110;
            15'b010010010010110 : data = 16'b0100111001011001;
            15'b010010010010111 : data = 16'b0100111001101100;
            15'b010010010011000 : data = 16'b0100111001111111;
            15'b010010010011001 : data = 16'b0100111010010010;
            15'b010010010011010 : data = 16'b0100111010100101;
            15'b010010010011011 : data = 16'b0100111010111000;
            15'b010010010011100 : data = 16'b0100111011001011;
            15'b010010010011101 : data = 16'b0100111011011110;
            15'b010010010011110 : data = 16'b0100111011110001;
            15'b010010010011111 : data = 16'b0100111100000100;
            15'b010010010100000 : data = 16'b0100111100010111;
            15'b010010010100001 : data = 16'b0100111100101010;
            15'b010010010100010 : data = 16'b0100111100111101;
            15'b010010010100011 : data = 16'b0100111101010000;
            15'b010010010100100 : data = 16'b0100111101100011;
            15'b010010010100101 : data = 16'b0100111101110110;
            15'b010010010100110 : data = 16'b0100111110001001;
            15'b010010010100111 : data = 16'b0100111110011100;
            15'b010010010101000 : data = 16'b0100111110101111;
            15'b010010010101001 : data = 16'b0100111111000011;
            15'b010010010101010 : data = 16'b0100111111010110;
            15'b010010010101011 : data = 16'b0100111111101001;
            15'b010010010101100 : data = 16'b0100111111111100;
            15'b010010010101101 : data = 16'b0101000000001111;
            15'b010010010101110 : data = 16'b0101000000100010;
            15'b010010010101111 : data = 16'b0101000000110101;
            15'b010010010110000 : data = 16'b0101000001001000;
            15'b010010010110001 : data = 16'b0101000001011011;
            15'b010010010110010 : data = 16'b0101000001101110;
            15'b010010010110011 : data = 16'b0101000010000010;
            15'b010010010110100 : data = 16'b0101000010010101;
            15'b010010010110101 : data = 16'b0101000010101000;
            15'b010010010110110 : data = 16'b0101000010111011;
            15'b010010010110111 : data = 16'b0101000011001110;
            15'b010010010111000 : data = 16'b0101000011100001;
            15'b010010010111001 : data = 16'b0101000011110100;
            15'b010010010111010 : data = 16'b0101000100000111;
            15'b010010010111011 : data = 16'b0101000100011011;
            15'b010010010111100 : data = 16'b0101000100101110;
            15'b010010010111101 : data = 16'b0101000101000001;
            15'b010010010111110 : data = 16'b0101000101010100;
            15'b010010010111111 : data = 16'b0101000101100111;
            15'b010010011000000 : data = 16'b0101000101111010;
            15'b010010011000001 : data = 16'b0101000110001110;
            15'b010010011000010 : data = 16'b0101000110100001;
            15'b010010011000011 : data = 16'b0101000110110100;
            15'b010010011000100 : data = 16'b0101000111000111;
            15'b010010011000101 : data = 16'b0101000111011010;
            15'b010010011000110 : data = 16'b0101000111101110;
            15'b010010011000111 : data = 16'b0101001000000001;
            15'b010010011001000 : data = 16'b0101001000010100;
            15'b010010011001001 : data = 16'b0101001000100111;
            15'b010010011001010 : data = 16'b0101001000111010;
            15'b010010011001011 : data = 16'b0101001001001110;
            15'b010010011001100 : data = 16'b0101001001100001;
            15'b010010011001101 : data = 16'b0101001001110100;
            15'b010010011001110 : data = 16'b0101001010000111;
            15'b010010011001111 : data = 16'b0101001010011011;
            15'b010010011010000 : data = 16'b0101001010101110;
            15'b010010011010001 : data = 16'b0101001011000001;
            15'b010010011010010 : data = 16'b0101001011010100;
            15'b010010011010011 : data = 16'b0101001011101000;
            15'b010010011010100 : data = 16'b0101001011111011;
            15'b010010011010101 : data = 16'b0101001100001110;
            15'b010010011010110 : data = 16'b0101001100100010;
            15'b010010011010111 : data = 16'b0101001100110101;
            15'b010010011011000 : data = 16'b0101001101001000;
            15'b010010011011001 : data = 16'b0101001101011011;
            15'b010010011011010 : data = 16'b0101001101101111;
            15'b010010011011011 : data = 16'b0101001110000010;
            15'b010010011011100 : data = 16'b0101001110010101;
            15'b010010011011101 : data = 16'b0101001110101001;
            15'b010010011011110 : data = 16'b0101001110111100;
            15'b010010011011111 : data = 16'b0101001111001111;
            15'b010010011100000 : data = 16'b0101001111100011;
            15'b010010011100001 : data = 16'b0101001111110110;
            15'b010010011100010 : data = 16'b0101010000001001;
            15'b010010011100011 : data = 16'b0101010000011101;
            15'b010010011100100 : data = 16'b0101010000110000;
            15'b010010011100101 : data = 16'b0101010001000011;
            15'b010010011100110 : data = 16'b0101010001010111;
            15'b010010011100111 : data = 16'b0101010001101010;
            15'b010010011101000 : data = 16'b0101010001111101;
            15'b010010011101001 : data = 16'b0101010010010001;
            15'b010010011101010 : data = 16'b0101010010100100;
            15'b010010011101011 : data = 16'b0101010010110111;
            15'b010010011101100 : data = 16'b0101010011001011;
            15'b010010011101101 : data = 16'b0101010011011110;
            15'b010010011101110 : data = 16'b0101010011110010;
            15'b010010011101111 : data = 16'b0101010100000101;
            15'b010010011110000 : data = 16'b0101010100011000;
            15'b010010011110001 : data = 16'b0101010100101100;
            15'b010010011110010 : data = 16'b0101010100111111;
            15'b010010011110011 : data = 16'b0101010101010011;
            15'b010010011110100 : data = 16'b0101010101100110;
            15'b010010011110101 : data = 16'b0101010101111001;
            15'b010010011110110 : data = 16'b0101010110001101;
            15'b010010011110111 : data = 16'b0101010110100000;
            15'b010010011111000 : data = 16'b0101010110110100;
            15'b010010011111001 : data = 16'b0101010111000111;
            15'b010010011111010 : data = 16'b0101010111011011;
            15'b010010011111011 : data = 16'b0101010111101110;
            15'b010010011111100 : data = 16'b0101011000000001;
            15'b010010011111101 : data = 16'b0101011000010101;
            15'b010010011111110 : data = 16'b0101011000101000;
            15'b010010011111111 : data = 16'b0101011000111100;
            15'b010010100000000 : data = 16'b0101011001001111;
            15'b010010100000001 : data = 16'b0101011001100011;
            15'b010010100000010 : data = 16'b0101011001110110;
            15'b010010100000011 : data = 16'b0101011010001010;
            15'b010010100000100 : data = 16'b0101011010011101;
            15'b010010100000101 : data = 16'b0101011010110001;
            15'b010010100000110 : data = 16'b0101011011000100;
            15'b010010100000111 : data = 16'b0101011011011000;
            15'b010010100001000 : data = 16'b0101011011101011;
            15'b010010100001001 : data = 16'b0101011011111111;
            15'b010010100001010 : data = 16'b0101011100010010;
            15'b010010100001011 : data = 16'b0101011100100110;
            15'b010010100001100 : data = 16'b0101011100111001;
            15'b010010100001101 : data = 16'b0101011101001101;
            15'b010010100001110 : data = 16'b0101011101100000;
            15'b010010100001111 : data = 16'b0101011101110100;
            15'b010010100010000 : data = 16'b0101011110000111;
            15'b010010100010001 : data = 16'b0101011110011011;
            15'b010010100010010 : data = 16'b0101011110101110;
            15'b010010100010011 : data = 16'b0101011111000010;
            15'b010010100010100 : data = 16'b0101011111010101;
            15'b010010100010101 : data = 16'b0101011111101001;
            15'b010010100010110 : data = 16'b0101011111111101;
            15'b010010100010111 : data = 16'b0101100000010000;
            15'b010010100011000 : data = 16'b0101100000100100;
            15'b010010100011001 : data = 16'b0101100000110111;
            15'b010010100011010 : data = 16'b0101100001001011;
            15'b010010100011011 : data = 16'b0101100001011110;
            15'b010010100011100 : data = 16'b0101100001110010;
            15'b010010100011101 : data = 16'b0101100010000110;
            15'b010010100011110 : data = 16'b0101100010011001;
            15'b010010100011111 : data = 16'b0101100010101101;
            15'b010010100100000 : data = 16'b0101100011000000;
            15'b010010100100001 : data = 16'b0101100011010100;
            15'b010010100100010 : data = 16'b0101100011100111;
            15'b010010100100011 : data = 16'b0101100011111011;
            15'b010010100100100 : data = 16'b0101100100001111;
            15'b010010100100101 : data = 16'b0101100100100010;
            15'b010010100100110 : data = 16'b0101100100110110;
            15'b010010100100111 : data = 16'b0101100101001010;
            15'b010010100101000 : data = 16'b0101100101011101;
            15'b010010100101001 : data = 16'b0101100101110001;
            15'b010010100101010 : data = 16'b0101100110000100;
            15'b010010100101011 : data = 16'b0101100110011000;
            15'b010010100101100 : data = 16'b0101100110101100;
            15'b010010100101101 : data = 16'b0101100110111111;
            15'b010010100101110 : data = 16'b0101100111010011;
            15'b010010100101111 : data = 16'b0101100111100111;
            15'b010010100110000 : data = 16'b0101100111111010;
            15'b010010100110001 : data = 16'b0101101000001110;
            15'b010010100110010 : data = 16'b0101101000100010;
            15'b010010100110011 : data = 16'b0101101000110101;
            15'b010010100110100 : data = 16'b0101101001001001;
            15'b010010100110101 : data = 16'b0101101001011101;
            15'b010010100110110 : data = 16'b0101101001110000;
            15'b010010100110111 : data = 16'b0101101010000100;
            15'b010010100111000 : data = 16'b0101101010011000;
            15'b010010100111001 : data = 16'b0101101010101011;
            15'b010010100111010 : data = 16'b0101101010111111;
            15'b010010100111011 : data = 16'b0101101011010011;
            15'b010010100111100 : data = 16'b0101101011100111;
            15'b010010100111101 : data = 16'b0101101011111010;
            15'b010010100111110 : data = 16'b0101101100001110;
            15'b010010100111111 : data = 16'b0101101100100010;
            15'b010010101000000 : data = 16'b0101101100110101;
            15'b010010101000001 : data = 16'b0101101101001001;
            15'b010010101000010 : data = 16'b0101101101011101;
            15'b010010101000011 : data = 16'b0101101101110001;
            15'b010010101000100 : data = 16'b0101101110000100;
            15'b010010101000101 : data = 16'b0101101110011000;
            15'b010010101000110 : data = 16'b0101101110101100;
            15'b010010101000111 : data = 16'b0101101110111111;
            15'b010010101001000 : data = 16'b0101101111010011;
            15'b010010101001001 : data = 16'b0101101111100111;
            15'b010010101001010 : data = 16'b0101101111111011;
            15'b010010101001011 : data = 16'b0101110000001111;
            15'b010010101001100 : data = 16'b0101110000100010;
            15'b010010101001101 : data = 16'b0101110000110110;
            15'b010010101001110 : data = 16'b0101110001001010;
            15'b010010101001111 : data = 16'b0101110001011110;
            15'b010010101010000 : data = 16'b0101110001110001;
            15'b010010101010001 : data = 16'b0101110010000101;
            15'b010010101010010 : data = 16'b0101110010011001;
            15'b010010101010011 : data = 16'b0101110010101101;
            15'b010010101010100 : data = 16'b0101110011000000;
            15'b010010101010101 : data = 16'b0101110011010100;
            15'b010010101010110 : data = 16'b0101110011101000;
            15'b010010101010111 : data = 16'b0101110011111100;
            15'b010010101011000 : data = 16'b0101110100010000;
            15'b010010101011001 : data = 16'b0101110100100011;
            15'b010010101011010 : data = 16'b0101110100110111;
            15'b010010101011011 : data = 16'b0101110101001011;
            15'b010010101011100 : data = 16'b0101110101011111;
            15'b010010101011101 : data = 16'b0101110101110011;
            15'b010010101011110 : data = 16'b0101110110000111;
            15'b010010101011111 : data = 16'b0101110110011010;
            15'b010010101100000 : data = 16'b0101110110101110;
            15'b010010101100001 : data = 16'b0101110111000010;
            15'b010010101100010 : data = 16'b0101110111010110;
            15'b010010101100011 : data = 16'b0101110111101010;
            15'b010010101100100 : data = 16'b0101110111111110;
            15'b010010101100101 : data = 16'b0101111000010001;
            15'b010010101100110 : data = 16'b0101111000100101;
            15'b010010101100111 : data = 16'b0101111000111001;
            15'b010010101101000 : data = 16'b0101111001001101;
            15'b010010101101001 : data = 16'b0101111001100001;
            15'b010010101101010 : data = 16'b0101111001110101;
            15'b010010101101011 : data = 16'b0101111010001001;
            15'b010010101101100 : data = 16'b0101111010011101;
            15'b010010101101101 : data = 16'b0101111010110000;
            15'b010010101101110 : data = 16'b0101111011000100;
            15'b010010101101111 : data = 16'b0101111011011000;
            15'b010010101110000 : data = 16'b0101111011101100;
            15'b010010101110001 : data = 16'b0101111100000000;
            15'b010010101110010 : data = 16'b0101111100010100;
            15'b010010101110011 : data = 16'b0101111100101000;
            15'b010010101110100 : data = 16'b0101111100111100;
            15'b010010101110101 : data = 16'b0101111101010000;
            15'b010010101110110 : data = 16'b0101111101100011;
            15'b010010101110111 : data = 16'b0101111101110111;
            15'b010010101111000 : data = 16'b0101111110001011;
            15'b010010101111001 : data = 16'b0101111110011111;
            15'b010010101111010 : data = 16'b0101111110110011;
            15'b010010101111011 : data = 16'b0101111111000111;
            15'b010010101111100 : data = 16'b0101111111011011;
            15'b010010101111101 : data = 16'b0101111111101111;
            15'b010010101111110 : data = 16'b0110000000000011;
            15'b010010101111111 : data = 16'b0110000000010111;
            15'b010010110000000 : data = 16'b0110000000101011;
            15'b010010110000001 : data = 16'b0110000000111111;
            15'b010010110000010 : data = 16'b0110000001010011;
            15'b010010110000011 : data = 16'b0110000001100111;
            15'b010010110000100 : data = 16'b0110000001111010;
            15'b010010110000101 : data = 16'b0110000010001110;
            15'b010010110000110 : data = 16'b0110000010100010;
            15'b010010110000111 : data = 16'b0110000010110110;
            15'b010010110001000 : data = 16'b0110000011001010;
            15'b010010110001001 : data = 16'b0110000011011110;
            15'b010010110001010 : data = 16'b0110000011110010;
            15'b010010110001011 : data = 16'b0110000100000110;
            15'b010010110001100 : data = 16'b0110000100011010;
            15'b010010110001101 : data = 16'b0110000100101110;
            15'b010010110001110 : data = 16'b0110000101000010;
            15'b010010110001111 : data = 16'b0110000101010110;
            15'b010010110010000 : data = 16'b0110000101101010;
            15'b010010110010001 : data = 16'b0110000101111110;
            15'b010010110010010 : data = 16'b0110000110010010;
            15'b010010110010011 : data = 16'b0110000110100110;
            15'b010010110010100 : data = 16'b0110000110111010;
            15'b010010110010101 : data = 16'b0110000111001110;
            15'b010010110010110 : data = 16'b0110000111100010;
            15'b010010110010111 : data = 16'b0110000111110110;
            15'b010010110011000 : data = 16'b0110001000001010;
            15'b010010110011001 : data = 16'b0110001000011110;
            15'b010010110011010 : data = 16'b0110001000110010;
            15'b010010110011011 : data = 16'b0110001001000110;
            15'b010010110011100 : data = 16'b0110001001011010;
            15'b010010110011101 : data = 16'b0110001001101110;
            15'b010010110011110 : data = 16'b0110001010000010;
            15'b010010110011111 : data = 16'b0110001010010110;
            15'b010010110100000 : data = 16'b0110001010101010;
            15'b010010110100001 : data = 16'b0110001010111110;
            15'b010010110100010 : data = 16'b0110001011010010;
            15'b010010110100011 : data = 16'b0110001011100111;
            15'b010010110100100 : data = 16'b0110001011111011;
            15'b010010110100101 : data = 16'b0110001100001111;
            15'b010010110100110 : data = 16'b0110001100100011;
            15'b010010110100111 : data = 16'b0110001100110111;
            15'b010010110101000 : data = 16'b0110001101001011;
            15'b010010110101001 : data = 16'b0110001101011111;
            15'b010010110101010 : data = 16'b0110001101110011;
            15'b010010110101011 : data = 16'b0110001110000111;
            15'b010010110101100 : data = 16'b0110001110011011;
            15'b010010110101101 : data = 16'b0110001110101111;
            15'b010010110101110 : data = 16'b0110001111000011;
            15'b010010110101111 : data = 16'b0110001111010111;
            15'b010010110110000 : data = 16'b0110001111101011;
            15'b010010110110001 : data = 16'b0110010000000000;
            15'b010010110110010 : data = 16'b0110010000010100;
            15'b010010110110011 : data = 16'b0110010000101000;
            15'b010010110110100 : data = 16'b0110010000111100;
            15'b010010110110101 : data = 16'b0110010001010000;
            15'b010010110110110 : data = 16'b0110010001100100;
            15'b010010110110111 : data = 16'b0110010001111000;
            15'b010010110111000 : data = 16'b0110010010001100;
            15'b010010110111001 : data = 16'b0110010010100000;
            15'b010010110111010 : data = 16'b0110010010110100;
            15'b010010110111011 : data = 16'b0110010011001001;
            15'b010010110111100 : data = 16'b0110010011011101;
            15'b010010110111101 : data = 16'b0110010011110001;
            15'b010010110111110 : data = 16'b0110010100000101;
            15'b010010110111111 : data = 16'b0110010100011001;
            15'b010010111000000 : data = 16'b0110010100101101;
            15'b010010111000001 : data = 16'b0110010101000001;
            15'b010010111000010 : data = 16'b0110010101010101;
            15'b010010111000011 : data = 16'b0110010101101010;
            15'b010010111000100 : data = 16'b0110010101111110;
            15'b010010111000101 : data = 16'b0110010110010010;
            15'b010010111000110 : data = 16'b0110010110100110;
            15'b010010111000111 : data = 16'b0110010110111010;
            15'b010010111001000 : data = 16'b0110010111001110;
            15'b010010111001001 : data = 16'b0110010111100010;
            15'b010010111001010 : data = 16'b0110010111110111;
            15'b010010111001011 : data = 16'b0110011000001011;
            15'b010010111001100 : data = 16'b0110011000011111;
            15'b010010111001101 : data = 16'b0110011000110011;
            15'b010010111001110 : data = 16'b0110011001000111;
            15'b010010111001111 : data = 16'b0110011001011011;
            15'b010010111010000 : data = 16'b0110011001110000;
            15'b010010111010001 : data = 16'b0110011010000100;
            15'b010010111010010 : data = 16'b0110011010011000;
            15'b010010111010011 : data = 16'b0110011010101100;
            15'b010010111010100 : data = 16'b0110011011000000;
            15'b010010111010101 : data = 16'b0110011011010101;
            15'b010010111010110 : data = 16'b0110011011101001;
            15'b010010111010111 : data = 16'b0110011011111101;
            15'b010010111011000 : data = 16'b0110011100010001;
            15'b010010111011001 : data = 16'b0110011100100101;
            15'b010010111011010 : data = 16'b0110011100111001;
            15'b010010111011011 : data = 16'b0110011101001110;
            15'b010010111011100 : data = 16'b0110011101100010;
            15'b010010111011101 : data = 16'b0110011101110110;
            15'b010010111011110 : data = 16'b0110011110001010;
            15'b010010111011111 : data = 16'b0110011110011110;
            15'b010010111100000 : data = 16'b0110011110110011;
            15'b010010111100001 : data = 16'b0110011111000111;
            15'b010010111100010 : data = 16'b0110011111011011;
            15'b010010111100011 : data = 16'b0110011111101111;
            15'b010010111100100 : data = 16'b0110100000000100;
            15'b010010111100101 : data = 16'b0110100000011000;
            15'b010010111100110 : data = 16'b0110100000101100;
            15'b010010111100111 : data = 16'b0110100001000000;
            15'b010010111101000 : data = 16'b0110100001010100;
            15'b010010111101001 : data = 16'b0110100001101001;
            15'b010010111101010 : data = 16'b0110100001111101;
            15'b010010111101011 : data = 16'b0110100010010001;
            15'b010010111101100 : data = 16'b0110100010100101;
            15'b010010111101101 : data = 16'b0110100010111010;
            15'b010010111101110 : data = 16'b0110100011001110;
            15'b010010111101111 : data = 16'b0110100011100010;
            15'b010010111110000 : data = 16'b0110100011110110;
            15'b010010111110001 : data = 16'b0110100100001011;
            15'b010010111110010 : data = 16'b0110100100011111;
            15'b010010111110011 : data = 16'b0110100100110011;
            15'b010010111110100 : data = 16'b0110100101000111;
            15'b010010111110101 : data = 16'b0110100101011100;
            15'b010010111110110 : data = 16'b0110100101110000;
            15'b010010111110111 : data = 16'b0110100110000100;
            15'b010010111111000 : data = 16'b0110100110011001;
            15'b010010111111001 : data = 16'b0110100110101101;
            15'b010010111111010 : data = 16'b0110100111000001;
            15'b010010111111011 : data = 16'b0110100111010101;
            15'b010010111111100 : data = 16'b0110100111101010;
            15'b010010111111101 : data = 16'b0110100111111110;
            15'b010010111111110 : data = 16'b0110101000010010;
            15'b010010111111111 : data = 16'b0110101000100110;
            15'b010011000000000 : data = 16'b0110101000111011;
            15'b010011000000001 : data = 16'b0110101001001111;
            15'b010011000000010 : data = 16'b0110101001100011;
            15'b010011000000011 : data = 16'b0110101001111000;
            15'b010011000000100 : data = 16'b0110101010001100;
            15'b010011000000101 : data = 16'b0110101010100000;
            15'b010011000000110 : data = 16'b0110101010110101;
            15'b010011000000111 : data = 16'b0110101011001001;
            15'b010011000001000 : data = 16'b0110101011011101;
            15'b010011000001001 : data = 16'b0110101011110001;
            15'b010011000001010 : data = 16'b0110101100000110;
            15'b010011000001011 : data = 16'b0110101100011010;
            15'b010011000001100 : data = 16'b0110101100101110;
            15'b010011000001101 : data = 16'b0110101101000011;
            15'b010011000001110 : data = 16'b0110101101010111;
            15'b010011000001111 : data = 16'b0110101101101011;
            15'b010011000010000 : data = 16'b0110101110000000;
            15'b010011000010001 : data = 16'b0110101110010100;
            15'b010011000010010 : data = 16'b0110101110101000;
            15'b010011000010011 : data = 16'b0110101110111101;
            15'b010011000010100 : data = 16'b0110101111010001;
            15'b010011000010101 : data = 16'b0110101111100101;
            15'b010011000010110 : data = 16'b0110101111111010;
            15'b010011000010111 : data = 16'b0110110000001110;
            15'b010011000011000 : data = 16'b0110110000100010;
            15'b010011000011001 : data = 16'b0110110000110111;
            15'b010011000011010 : data = 16'b0110110001001011;
            15'b010011000011011 : data = 16'b0110110001011111;
            15'b010011000011100 : data = 16'b0110110001110100;
            15'b010011000011101 : data = 16'b0110110010001000;
            15'b010011000011110 : data = 16'b0110110010011100;
            15'b010011000011111 : data = 16'b0110110010110001;
            15'b010011000100000 : data = 16'b0110110011000101;
            15'b010011000100001 : data = 16'b0110110011011001;
            15'b010011000100010 : data = 16'b0110110011101110;
            15'b010011000100011 : data = 16'b0110110100000010;
            15'b010011000100100 : data = 16'b0110110100010110;
            15'b010011000100101 : data = 16'b0110110100101011;
            15'b010011000100110 : data = 16'b0110110100111111;
            15'b010011000100111 : data = 16'b0110110101010100;
            15'b010011000101000 : data = 16'b0110110101101000;
            15'b010011000101001 : data = 16'b0110110101111100;
            15'b010011000101010 : data = 16'b0110110110010001;
            15'b010011000101011 : data = 16'b0110110110100101;
            15'b010011000101100 : data = 16'b0110110110111001;
            15'b010011000101101 : data = 16'b0110110111001110;
            15'b010011000101110 : data = 16'b0110110111100010;
            15'b010011000101111 : data = 16'b0110110111110111;
            15'b010011000110000 : data = 16'b0110111000001011;
            15'b010011000110001 : data = 16'b0110111000011111;
            15'b010011000110010 : data = 16'b0110111000110100;
            15'b010011000110011 : data = 16'b0110111001001000;
            15'b010011000110100 : data = 16'b0110111001011101;
            15'b010011000110101 : data = 16'b0110111001110001;
            15'b010011000110110 : data = 16'b0110111010000101;
            15'b010011000110111 : data = 16'b0110111010011010;
            15'b010011000111000 : data = 16'b0110111010101110;
            15'b010011000111001 : data = 16'b0110111011000011;
            15'b010011000111010 : data = 16'b0110111011010111;
            15'b010011000111011 : data = 16'b0110111011101011;
            15'b010011000111100 : data = 16'b0110111100000000;
            15'b010011000111101 : data = 16'b0110111100010100;
            15'b010011000111110 : data = 16'b0110111100101001;
            15'b010011000111111 : data = 16'b0110111100111101;
            15'b010011001000000 : data = 16'b0110111101010001;
            15'b010011001000001 : data = 16'b0110111101100110;
            15'b010011001000010 : data = 16'b0110111101111010;
            15'b010011001000011 : data = 16'b0110111110001111;
            15'b010011001000100 : data = 16'b0110111110100011;
            15'b010011001000101 : data = 16'b0110111110110111;
            15'b010011001000110 : data = 16'b0110111111001100;
            15'b010011001000111 : data = 16'b0110111111100000;
            15'b010011001001000 : data = 16'b0110111111110101;
            15'b010011001001001 : data = 16'b0111000000001001;
            15'b010011001001010 : data = 16'b0111000000011110;
            15'b010011001001011 : data = 16'b0111000000110010;
            15'b010011001001100 : data = 16'b0111000001000110;
            15'b010011001001101 : data = 16'b0111000001011011;
            15'b010011001001110 : data = 16'b0111000001101111;
            15'b010011001001111 : data = 16'b0111000010000100;
            15'b010011001010000 : data = 16'b0111000010011000;
            15'b010011001010001 : data = 16'b0111000010101101;
            15'b010011001010010 : data = 16'b0111000011000001;
            15'b010011001010011 : data = 16'b0111000011010101;
            15'b010011001010100 : data = 16'b0111000011101010;
            15'b010011001010101 : data = 16'b0111000011111110;
            15'b010011001010110 : data = 16'b0111000100010011;
            15'b010011001010111 : data = 16'b0111000100100111;
            15'b010011001011000 : data = 16'b0111000100111100;
            15'b010011001011001 : data = 16'b0111000101010000;
            15'b010011001011010 : data = 16'b0111000101100101;
            15'b010011001011011 : data = 16'b0111000101111001;
            15'b010011001011100 : data = 16'b0111000110001110;
            15'b010011001011101 : data = 16'b0111000110100010;
            15'b010011001011110 : data = 16'b0111000110110110;
            15'b010011001011111 : data = 16'b0111000111001011;
            15'b010011001100000 : data = 16'b0111000111011111;
            15'b010011001100001 : data = 16'b0111000111110100;
            15'b010011001100010 : data = 16'b0111001000001000;
            15'b010011001100011 : data = 16'b0111001000011101;
            15'b010011001100100 : data = 16'b0111001000110001;
            15'b010011001100101 : data = 16'b0111001001000110;
            15'b010011001100110 : data = 16'b0111001001011010;
            15'b010011001100111 : data = 16'b0111001001101111;
            15'b010011001101000 : data = 16'b0111001010000011;
            15'b010011001101001 : data = 16'b0111001010011000;
            15'b010011001101010 : data = 16'b0111001010101100;
            15'b010011001101011 : data = 16'b0111001011000001;
            15'b010011001101100 : data = 16'b0111001011010101;
            15'b010011001101101 : data = 16'b0111001011101010;
            15'b010011001101110 : data = 16'b0111001011111110;
            15'b010011001101111 : data = 16'b0111001100010010;
            15'b010011001110000 : data = 16'b0111001100100111;
            15'b010011001110001 : data = 16'b0111001100111011;
            15'b010011001110010 : data = 16'b0111001101010000;
            15'b010011001110011 : data = 16'b0111001101100100;
            15'b010011001110100 : data = 16'b0111001101111001;
            15'b010011001110101 : data = 16'b0111001110001101;
            15'b010011001110110 : data = 16'b0111001110100010;
            15'b010011001110111 : data = 16'b0111001110110110;
            15'b010011001111000 : data = 16'b0111001111001011;
            15'b010011001111001 : data = 16'b0111001111011111;
            15'b010011001111010 : data = 16'b0111001111110100;
            15'b010011001111011 : data = 16'b0111010000001000;
            15'b010011001111100 : data = 16'b0111010000011101;
            15'b010011001111101 : data = 16'b0111010000110001;
            15'b010011001111110 : data = 16'b0111010001000110;
            15'b010011001111111 : data = 16'b0111010001011010;
            15'b010011010000000 : data = 16'b0111010001101111;
            15'b010011010000001 : data = 16'b0111010010000011;
            15'b010011010000010 : data = 16'b0111010010011000;
            15'b010011010000011 : data = 16'b0111010010101100;
            15'b010011010000100 : data = 16'b0111010011000001;
            15'b010011010000101 : data = 16'b0111010011010101;
            15'b010011010000110 : data = 16'b0111010011101010;
            15'b010011010000111 : data = 16'b0111010011111110;
            15'b010011010001000 : data = 16'b0111010100010011;
            15'b010011010001001 : data = 16'b0111010100100111;
            15'b010011010001010 : data = 16'b0111010100111100;
            15'b010011010001011 : data = 16'b0111010101010000;
            15'b010011010001100 : data = 16'b0111010101100101;
            15'b010011010001101 : data = 16'b0111010101111010;
            15'b010011010001110 : data = 16'b0111010110001110;
            15'b010011010001111 : data = 16'b0111010110100011;
            15'b010011010010000 : data = 16'b0111010110110111;
            15'b010011010010001 : data = 16'b0111010111001100;
            15'b010011010010010 : data = 16'b0111010111100000;
            15'b010011010010011 : data = 16'b0111010111110101;
            15'b010011010010100 : data = 16'b0111011000001001;
            15'b010011010010101 : data = 16'b0111011000011110;
            15'b010011010010110 : data = 16'b0111011000110010;
            15'b010011010010111 : data = 16'b0111011001000111;
            15'b010011010011000 : data = 16'b0111011001011011;
            15'b010011010011001 : data = 16'b0111011001110000;
            15'b010011010011010 : data = 16'b0111011010000100;
            15'b010011010011011 : data = 16'b0111011010011001;
            15'b010011010011100 : data = 16'b0111011010101101;
            15'b010011010011101 : data = 16'b0111011011000010;
            15'b010011010011110 : data = 16'b0111011011010110;
            15'b010011010011111 : data = 16'b0111011011101011;
            15'b010011010100000 : data = 16'b0111011100000000;
            15'b010011010100001 : data = 16'b0111011100010100;
            15'b010011010100010 : data = 16'b0111011100101001;
            15'b010011010100011 : data = 16'b0111011100111101;
            15'b010011010100100 : data = 16'b0111011101010010;
            15'b010011010100101 : data = 16'b0111011101100110;
            15'b010011010100110 : data = 16'b0111011101111011;
            15'b010011010100111 : data = 16'b0111011110001111;
            15'b010011010101000 : data = 16'b0111011110100100;
            15'b010011010101001 : data = 16'b0111011110111000;
            15'b010011010101010 : data = 16'b0111011111001101;
            15'b010011010101011 : data = 16'b0111011111100001;
            15'b010011010101100 : data = 16'b0111011111110110;
            15'b010011010101101 : data = 16'b0111100000001011;
            15'b010011010101110 : data = 16'b0111100000011111;
            15'b010011010101111 : data = 16'b0111100000110100;
            15'b010011010110000 : data = 16'b0111100001001000;
            15'b010011010110001 : data = 16'b0111100001011101;
            15'b010011010110010 : data = 16'b0111100001110001;
            15'b010011010110011 : data = 16'b0111100010000110;
            15'b010011010110100 : data = 16'b0111100010011010;
            15'b010011010110101 : data = 16'b0111100010101111;
            15'b010011010110110 : data = 16'b0111100011000100;
            15'b010011010110111 : data = 16'b0111100011011000;
            15'b010011010111000 : data = 16'b0111100011101101;
            15'b010011010111001 : data = 16'b0111100100000001;
            15'b010011010111010 : data = 16'b0111100100010110;
            15'b010011010111011 : data = 16'b0111100100101010;
            15'b010011010111100 : data = 16'b0111100100111111;
            15'b010011010111101 : data = 16'b0111100101010011;
            15'b010011010111110 : data = 16'b0111100101101000;
            15'b010011010111111 : data = 16'b0111100101111101;
            15'b010011011000000 : data = 16'b0111100110010001;
            15'b010011011000001 : data = 16'b0111100110100110;
            15'b010011011000010 : data = 16'b0111100110111010;
            15'b010011011000011 : data = 16'b0111100111001111;
            15'b010011011000100 : data = 16'b0111100111100011;
            15'b010011011000101 : data = 16'b0111100111111000;
            15'b010011011000110 : data = 16'b0111101000001101;
            15'b010011011000111 : data = 16'b0111101000100001;
            15'b010011011001000 : data = 16'b0111101000110110;
            15'b010011011001001 : data = 16'b0111101001001010;
            15'b010011011001010 : data = 16'b0111101001011111;
            15'b010011011001011 : data = 16'b0111101001110011;
            15'b010011011001100 : data = 16'b0111101010001000;
            15'b010011011001101 : data = 16'b0111101010011101;
            15'b010011011001110 : data = 16'b0111101010110001;
            15'b010011011001111 : data = 16'b0111101011000110;
            15'b010011011010000 : data = 16'b0111101011011010;
            15'b010011011010001 : data = 16'b0111101011101111;
            15'b010011011010010 : data = 16'b0111101100000011;
            15'b010011011010011 : data = 16'b0111101100011000;
            15'b010011011010100 : data = 16'b0111101100101101;
            15'b010011011010101 : data = 16'b0111101101000001;
            15'b010011011010110 : data = 16'b0111101101010110;
            15'b010011011010111 : data = 16'b0111101101101010;
            15'b010011011011000 : data = 16'b0111101101111111;
            15'b010011011011001 : data = 16'b0111101110010011;
            15'b010011011011010 : data = 16'b0111101110101000;
            15'b010011011011011 : data = 16'b0111101110111101;
            15'b010011011011100 : data = 16'b0111101111010001;
            15'b010011011011101 : data = 16'b0111101111100110;
            15'b010011011011110 : data = 16'b0111101111111010;
            15'b010011011011111 : data = 16'b0111110000001111;
            15'b010011011100000 : data = 16'b0111110000100011;
            15'b010011011100001 : data = 16'b0111110000111000;
            15'b010011011100010 : data = 16'b0111110001001101;
            15'b010011011100011 : data = 16'b0111110001100001;
            15'b010011011100100 : data = 16'b0111110001110110;
            15'b010011011100101 : data = 16'b0111110010001010;
            15'b010011011100110 : data = 16'b0111110010011111;
            15'b010011011100111 : data = 16'b0111110010110011;
            15'b010011011101000 : data = 16'b0111110011001000;
            15'b010011011101001 : data = 16'b0111110011011101;
            15'b010011011101010 : data = 16'b0111110011110001;
            15'b010011011101011 : data = 16'b0111110100000110;
            15'b010011011101100 : data = 16'b0111110100011010;
            15'b010011011101101 : data = 16'b0111110100101111;
            15'b010011011101110 : data = 16'b0111110101000100;
            15'b010011011101111 : data = 16'b0111110101011000;
            15'b010011011110000 : data = 16'b0111110101101101;
            15'b010011011110001 : data = 16'b0111110110000001;
            15'b010011011110010 : data = 16'b0111110110010110;
            15'b010011011110011 : data = 16'b0111110110101010;
            15'b010011011110100 : data = 16'b0111110110111111;
            15'b010011011110101 : data = 16'b0111110111010100;
            15'b010011011110110 : data = 16'b0111110111101000;
            15'b010011011110111 : data = 16'b0111110111111101;
            15'b010011011111000 : data = 16'b0111111000010001;
            15'b010011011111001 : data = 16'b0111111000100110;
            15'b010011011111010 : data = 16'b0111111000111011;
            15'b010011011111011 : data = 16'b0111111001001111;
            15'b010011011111100 : data = 16'b0111111001100100;
            15'b010011011111101 : data = 16'b0111111001111000;
            15'b010011011111110 : data = 16'b0111111010001101;
            15'b010011011111111 : data = 16'b0111111010100010;
            15'b010011100000000 : data = 16'b0111111010110110;
            15'b010011100000001 : data = 16'b0111111011001011;
            15'b010011100000010 : data = 16'b0111111011011111;
            15'b010011100000011 : data = 16'b0111111011110100;
            15'b010011100000100 : data = 16'b0111111100001000;
            15'b010011100000101 : data = 16'b0111111100011101;
            15'b010011100000110 : data = 16'b0111111100110010;
            15'b010011100000111 : data = 16'b0111111101000110;
            15'b010011100001000 : data = 16'b0111111101011011;
            15'b010011100001001 : data = 16'b0111111101101111;
            15'b010011100001010 : data = 16'b0111111110000100;
            15'b010011100001011 : data = 16'b0111111110011001;
            15'b010011100001100 : data = 16'b0111111110101101;
            15'b010011100001101 : data = 16'b0111111111000010;
            15'b010011100001110 : data = 16'b0111111111010110;
            15'b010011100001111 : data = 16'b0111111111101011;
            default : data = 16'b0000000000000000;
        endcase
    end
endmodule
