module memory (
    input [13:0] addr1,
    input [13:0] addr2,
    input [13:0] addr3,
    output reg [11:0] data1,
    output reg [11:0] data2,
    output reg [11:0] data3
);

    reg [11:0] mem [0:9999];

    initial begin
        mem[0] = 12'b000000000000;
        mem[1] = 12'b000000000000;
        mem[2] = 12'b000000000001;
        mem[3] = 12'b000000000001;
        mem[4] = 12'b000000000010;
        mem[5] = 12'b000000000011;
        mem[6] = 12'b000000000011;
        mem[7] = 12'b000000000100;
        mem[8] = 12'b000000000101;
        mem[9] = 12'b000000000101;
        mem[10] = 12'b000000000110;
        mem[11] = 12'b000000000111;
        mem[12] = 12'b000000000111;
        mem[13] = 12'b000000001000;
        mem[14] = 12'b000000001001;
        mem[15] = 12'b000000001001;
        mem[16] = 12'b000000001010;
        mem[17] = 12'b000000001010;
        mem[18] = 12'b000000001011;
        mem[19] = 12'b000000001100;
        mem[20] = 12'b000000001100;
        mem[21] = 12'b000000001101;
        mem[22] = 12'b000000001110;
        mem[23] = 12'b000000001110;
        mem[24] = 12'b000000001111;
        mem[25] = 12'b000000010000;
        mem[26] = 12'b000000010000;
        mem[27] = 12'b000000010001;
        mem[28] = 12'b000000010010;
        mem[29] = 12'b000000010010;
        mem[30] = 12'b000000010011;
        mem[31] = 12'b000000010011;
        mem[32] = 12'b000000010100;
        mem[33] = 12'b000000010101;
        mem[34] = 12'b000000010101;
        mem[35] = 12'b000000010110;
        mem[36] = 12'b000000010111;
        mem[37] = 12'b000000010111;
        mem[38] = 12'b000000011000;
        mem[39] = 12'b000000011001;
        mem[40] = 12'b000000011001;
        mem[41] = 12'b000000011010;
        mem[42] = 12'b000000011011;
        mem[43] = 12'b000000011011;
        mem[44] = 12'b000000011100;
        mem[45] = 12'b000000011100;
        mem[46] = 12'b000000011101;
        mem[47] = 12'b000000011110;
        mem[48] = 12'b000000011110;
        mem[49] = 12'b000000011111;
        mem[50] = 12'b000000100000;
        mem[51] = 12'b000000100000;
        mem[52] = 12'b000000100001;
        mem[53] = 12'b000000100010;
        mem[54] = 12'b000000100010;
        mem[55] = 12'b000000100011;
        mem[56] = 12'b000000100100;
        mem[57] = 12'b000000100100;
        mem[58] = 12'b000000100101;
        mem[59] = 12'b000000100101;
        mem[60] = 12'b000000100110;
        mem[61] = 12'b000000100111;
        mem[62] = 12'b000000100111;
        mem[63] = 12'b000000101000;
        mem[64] = 12'b000000101001;
        mem[65] = 12'b000000101001;
        mem[66] = 12'b000000101010;
        mem[67] = 12'b000000101011;
        mem[68] = 12'b000000101011;
        mem[69] = 12'b000000101100;
        mem[70] = 12'b000000101101;
        mem[71] = 12'b000000101101;
        mem[72] = 12'b000000101110;
        mem[73] = 12'b000000101110;
        mem[74] = 12'b000000101111;
        mem[75] = 12'b000000110000;
        mem[76] = 12'b000000110000;
        mem[77] = 12'b000000110001;
        mem[78] = 12'b000000110010;
        mem[79] = 12'b000000110010;
        mem[80] = 12'b000000110011;
        mem[81] = 12'b000000110100;
        mem[82] = 12'b000000110100;
        mem[83] = 12'b000000110101;
        mem[84] = 12'b000000110110;
        mem[85] = 12'b000000110110;
        mem[86] = 12'b000000110111;
        mem[87] = 12'b000000110111;
        mem[88] = 12'b000000111000;
        mem[89] = 12'b000000111001;
        mem[90] = 12'b000000111001;
        mem[91] = 12'b000000111010;
        mem[92] = 12'b000000111011;
        mem[93] = 12'b000000111011;
        mem[94] = 12'b000000111100;
        mem[95] = 12'b000000111101;
        mem[96] = 12'b000000111101;
        mem[97] = 12'b000000111110;
        mem[98] = 12'b000000111111;
        mem[99] = 12'b000000111111;
        mem[100] = 12'b000001000000;
        mem[101] = 12'b000001000000;
        mem[102] = 12'b000001000001;
        mem[103] = 12'b000001000010;
        mem[104] = 12'b000001000010;
        mem[105] = 12'b000001000011;
        mem[106] = 12'b000001000100;
        mem[107] = 12'b000001000100;
        mem[108] = 12'b000001000101;
        mem[109] = 12'b000001000110;
        mem[110] = 12'b000001000110;
        mem[111] = 12'b000001000111;
        mem[112] = 12'b000001001000;
        mem[113] = 12'b000001001000;
        mem[114] = 12'b000001001001;
        mem[115] = 12'b000001001001;
        mem[116] = 12'b000001001010;
        mem[117] = 12'b000001001011;
        mem[118] = 12'b000001001011;
        mem[119] = 12'b000001001100;
        mem[120] = 12'b000001001101;
        mem[121] = 12'b000001001101;
        mem[122] = 12'b000001001110;
        mem[123] = 12'b000001001111;
        mem[124] = 12'b000001001111;
        mem[125] = 12'b000001010000;
        mem[126] = 12'b000001010001;
        mem[127] = 12'b000001010001;
        mem[128] = 12'b000001010010;
        mem[129] = 12'b000001010010;
        mem[130] = 12'b000001010011;
        mem[131] = 12'b000001010100;
        mem[132] = 12'b000001010100;
        mem[133] = 12'b000001010101;
        mem[134] = 12'b000001010110;
        mem[135] = 12'b000001010110;
        mem[136] = 12'b000001010111;
        mem[137] = 12'b000001011000;
        mem[138] = 12'b000001011000;
        mem[139] = 12'b000001011001;
        mem[140] = 12'b000001011010;
        mem[141] = 12'b000001011010;
        mem[142] = 12'b000001011011;
        mem[143] = 12'b000001011011;
        mem[144] = 12'b000001011100;
        mem[145] = 12'b000001011101;
        mem[146] = 12'b000001011101;
        mem[147] = 12'b000001011110;
        mem[148] = 12'b000001011111;
        mem[149] = 12'b000001011111;
        mem[150] = 12'b000001100000;
        mem[151] = 12'b000001100001;
        mem[152] = 12'b000001100001;
        mem[153] = 12'b000001100010;
        mem[154] = 12'b000001100011;
        mem[155] = 12'b000001100011;
        mem[156] = 12'b000001100100;
        mem[157] = 12'b000001100100;
        mem[158] = 12'b000001100101;
        mem[159] = 12'b000001100110;
        mem[160] = 12'b000001100110;
        mem[161] = 12'b000001100111;
        mem[162] = 12'b000001101000;
        mem[163] = 12'b000001101000;
        mem[164] = 12'b000001101001;
        mem[165] = 12'b000001101010;
        mem[166] = 12'b000001101010;
        mem[167] = 12'b000001101011;
        mem[168] = 12'b000001101011;
        mem[169] = 12'b000001101100;
        mem[170] = 12'b000001101101;
        mem[171] = 12'b000001101101;
        mem[172] = 12'b000001101110;
        mem[173] = 12'b000001101111;
        mem[174] = 12'b000001101111;
        mem[175] = 12'b000001110000;
        mem[176] = 12'b000001110001;
        mem[177] = 12'b000001110001;
        mem[178] = 12'b000001110010;
        mem[179] = 12'b000001110011;
        mem[180] = 12'b000001110011;
        mem[181] = 12'b000001110100;
        mem[182] = 12'b000001110100;
        mem[183] = 12'b000001110101;
        mem[184] = 12'b000001110110;
        mem[185] = 12'b000001110110;
        mem[186] = 12'b000001110111;
        mem[187] = 12'b000001111000;
        mem[188] = 12'b000001111000;
        mem[189] = 12'b000001111001;
        mem[190] = 12'b000001111010;
        mem[191] = 12'b000001111010;
        mem[192] = 12'b000001111011;
        mem[193] = 12'b000001111100;
        mem[194] = 12'b000001111100;
        mem[195] = 12'b000001111101;
        mem[196] = 12'b000001111101;
        mem[197] = 12'b000001111110;
        mem[198] = 12'b000001111111;
        mem[199] = 12'b000001111111;
        mem[200] = 12'b000010000000;
        mem[201] = 12'b000010000001;
        mem[202] = 12'b000010000001;
        mem[203] = 12'b000010000010;
        mem[204] = 12'b000010000011;
        mem[205] = 12'b000010000011;
        mem[206] = 12'b000010000100;
        mem[207] = 12'b000010000101;
        mem[208] = 12'b000010000101;
        mem[209] = 12'b000010000110;
        mem[210] = 12'b000010000110;
        mem[211] = 12'b000010000111;
        mem[212] = 12'b000010001000;
        mem[213] = 12'b000010001000;
        mem[214] = 12'b000010001001;
        mem[215] = 12'b000010001010;
        mem[216] = 12'b000010001010;
        mem[217] = 12'b000010001011;
        mem[218] = 12'b000010001100;
        mem[219] = 12'b000010001100;
        mem[220] = 12'b000010001101;
        mem[221] = 12'b000010001110;
        mem[222] = 12'b000010001110;
        mem[223] = 12'b000010001111;
        mem[224] = 12'b000010001111;
        mem[225] = 12'b000010010000;
        mem[226] = 12'b000010010001;
        mem[227] = 12'b000010010001;
        mem[228] = 12'b000010010010;
        mem[229] = 12'b000010010011;
        mem[230] = 12'b000010010011;
        mem[231] = 12'b000010010100;
        mem[232] = 12'b000010010101;
        mem[233] = 12'b000010010101;
        mem[234] = 12'b000010010110;
        mem[235] = 12'b000010010111;
        mem[236] = 12'b000010010111;
        mem[237] = 12'b000010011000;
        mem[238] = 12'b000010011000;
        mem[239] = 12'b000010011001;
        mem[240] = 12'b000010011010;
        mem[241] = 12'b000010011010;
        mem[242] = 12'b000010011011;
        mem[243] = 12'b000010011100;
        mem[244] = 12'b000010011100;
        mem[245] = 12'b000010011101;
        mem[246] = 12'b000010011110;
        mem[247] = 12'b000010011110;
        mem[248] = 12'b000010011111;
        mem[249] = 12'b000010011111;
        mem[250] = 12'b000010100000;
        mem[251] = 12'b000010100001;
        mem[252] = 12'b000010100001;
        mem[253] = 12'b000010100010;
        mem[254] = 12'b000010100011;
        mem[255] = 12'b000010100011;
        mem[256] = 12'b000010100100;
        mem[257] = 12'b000010100101;
        mem[258] = 12'b000010100101;
        mem[259] = 12'b000010100110;
        mem[260] = 12'b000010100111;
        mem[261] = 12'b000010100111;
        mem[262] = 12'b000010101000;
        mem[263] = 12'b000010101000;
        mem[264] = 12'b000010101001;
        mem[265] = 12'b000010101010;
        mem[266] = 12'b000010101010;
        mem[267] = 12'b000010101011;
        mem[268] = 12'b000010101100;
        mem[269] = 12'b000010101100;
        mem[270] = 12'b000010101101;
        mem[271] = 12'b000010101110;
        mem[272] = 12'b000010101110;
        mem[273] = 12'b000010101111;
        mem[274] = 12'b000010110000;
        mem[275] = 12'b000010110000;
        mem[276] = 12'b000010110001;
        mem[277] = 12'b000010110001;
        mem[278] = 12'b000010110010;
        mem[279] = 12'b000010110011;
        mem[280] = 12'b000010110011;
        mem[281] = 12'b000010110100;
        mem[282] = 12'b000010110101;
        mem[283] = 12'b000010110101;
        mem[284] = 12'b000010110110;
        mem[285] = 12'b000010110111;
        mem[286] = 12'b000010110111;
        mem[287] = 12'b000010111000;
        mem[288] = 12'b000010111000;
        mem[289] = 12'b000010111001;
        mem[290] = 12'b000010111010;
        mem[291] = 12'b000010111010;
        mem[292] = 12'b000010111011;
        mem[293] = 12'b000010111100;
        mem[294] = 12'b000010111100;
        mem[295] = 12'b000010111101;
        mem[296] = 12'b000010111110;
        mem[297] = 12'b000010111110;
        mem[298] = 12'b000010111111;
        mem[299] = 12'b000011000000;
        mem[300] = 12'b000011000000;
        mem[301] = 12'b000011000001;
        mem[302] = 12'b000011000001;
        mem[303] = 12'b000011000010;
        mem[304] = 12'b000011000011;
        mem[305] = 12'b000011000011;
        mem[306] = 12'b000011000100;
        mem[307] = 12'b000011000101;
        mem[308] = 12'b000011000101;
        mem[309] = 12'b000011000110;
        mem[310] = 12'b000011000111;
        mem[311] = 12'b000011000111;
        mem[312] = 12'b000011001000;
        mem[313] = 12'b000011001000;
        mem[314] = 12'b000011001001;
        mem[315] = 12'b000011001010;
        mem[316] = 12'b000011001010;
        mem[317] = 12'b000011001011;
        mem[318] = 12'b000011001100;
        mem[319] = 12'b000011001100;
        mem[320] = 12'b000011001101;
        mem[321] = 12'b000011001110;
        mem[322] = 12'b000011001110;
        mem[323] = 12'b000011001111;
        mem[324] = 12'b000011010000;
        mem[325] = 12'b000011010000;
        mem[326] = 12'b000011010001;
        mem[327] = 12'b000011010001;
        mem[328] = 12'b000011010010;
        mem[329] = 12'b000011010011;
        mem[330] = 12'b000011010011;
        mem[331] = 12'b000011010100;
        mem[332] = 12'b000011010101;
        mem[333] = 12'b000011010101;
        mem[334] = 12'b000011010110;
        mem[335] = 12'b000011010111;
        mem[336] = 12'b000011010111;
        mem[337] = 12'b000011011000;
        mem[338] = 12'b000011011000;
        mem[339] = 12'b000011011001;
        mem[340] = 12'b000011011010;
        mem[341] = 12'b000011011010;
        mem[342] = 12'b000011011011;
        mem[343] = 12'b000011011100;
        mem[344] = 12'b000011011100;
        mem[345] = 12'b000011011101;
        mem[346] = 12'b000011011110;
        mem[347] = 12'b000011011110;
        mem[348] = 12'b000011011111;
        mem[349] = 12'b000011100000;
        mem[350] = 12'b000011100000;
        mem[351] = 12'b000011100001;
        mem[352] = 12'b000011100001;
        mem[353] = 12'b000011100010;
        mem[354] = 12'b000011100011;
        mem[355] = 12'b000011100011;
        mem[356] = 12'b000011100100;
        mem[357] = 12'b000011100101;
        mem[358] = 12'b000011100101;
        mem[359] = 12'b000011100110;
        mem[360] = 12'b000011100111;
        mem[361] = 12'b000011100111;
        mem[362] = 12'b000011101000;
        mem[363] = 12'b000011101000;
        mem[364] = 12'b000011101001;
        mem[365] = 12'b000011101010;
        mem[366] = 12'b000011101010;
        mem[367] = 12'b000011101011;
        mem[368] = 12'b000011101100;
        mem[369] = 12'b000011101100;
        mem[370] = 12'b000011101101;
        mem[371] = 12'b000011101110;
        mem[372] = 12'b000011101110;
        mem[373] = 12'b000011101111;
        mem[374] = 12'b000011101111;
        mem[375] = 12'b000011110000;
        mem[376] = 12'b000011110001;
        mem[377] = 12'b000011110001;
        mem[378] = 12'b000011110010;
        mem[379] = 12'b000011110011;
        mem[380] = 12'b000011110011;
        mem[381] = 12'b000011110100;
        mem[382] = 12'b000011110101;
        mem[383] = 12'b000011110101;
        mem[384] = 12'b000011110110;
        mem[385] = 12'b000011110111;
        mem[386] = 12'b000011110111;
        mem[387] = 12'b000011111000;
        mem[388] = 12'b000011111000;
        mem[389] = 12'b000011111001;
        mem[390] = 12'b000011111010;
        mem[391] = 12'b000011111010;
        mem[392] = 12'b000011111011;
        mem[393] = 12'b000011111100;
        mem[394] = 12'b000011111100;
        mem[395] = 12'b000011111101;
        mem[396] = 12'b000011111110;
        mem[397] = 12'b000011111110;
        mem[398] = 12'b000011111111;
        mem[399] = 12'b000011111111;
        mem[400] = 12'b000100000000;
        mem[401] = 12'b000100000001;
        mem[402] = 12'b000100000001;
        mem[403] = 12'b000100000010;
        mem[404] = 12'b000100000011;
        mem[405] = 12'b000100000011;
        mem[406] = 12'b000100000100;
        mem[407] = 12'b000100000101;
        mem[408] = 12'b000100000101;
        mem[409] = 12'b000100000110;
        mem[410] = 12'b000100000110;
        mem[411] = 12'b000100000111;
        mem[412] = 12'b000100001000;
        mem[413] = 12'b000100001000;
        mem[414] = 12'b000100001001;
        mem[415] = 12'b000100001010;
        mem[416] = 12'b000100001010;
        mem[417] = 12'b000100001011;
        mem[418] = 12'b000100001100;
        mem[419] = 12'b000100001100;
        mem[420] = 12'b000100001101;
        mem[421] = 12'b000100001101;
        mem[422] = 12'b000100001110;
        mem[423] = 12'b000100001111;
        mem[424] = 12'b000100001111;
        mem[425] = 12'b000100010000;
        mem[426] = 12'b000100010001;
        mem[427] = 12'b000100010001;
        mem[428] = 12'b000100010010;
        mem[429] = 12'b000100010011;
        mem[430] = 12'b000100010011;
        mem[431] = 12'b000100010100;
        mem[432] = 12'b000100010100;
        mem[433] = 12'b000100010101;
        mem[434] = 12'b000100010110;
        mem[435] = 12'b000100010110;
        mem[436] = 12'b000100010111;
        mem[437] = 12'b000100011000;
        mem[438] = 12'b000100011000;
        mem[439] = 12'b000100011001;
        mem[440] = 12'b000100011010;
        mem[441] = 12'b000100011010;
        mem[442] = 12'b000100011011;
        mem[443] = 12'b000100011011;
        mem[444] = 12'b000100011100;
        mem[445] = 12'b000100011101;
        mem[446] = 12'b000100011101;
        mem[447] = 12'b000100011110;
        mem[448] = 12'b000100011111;
        mem[449] = 12'b000100011111;
        mem[450] = 12'b000100100000;
        mem[451] = 12'b000100100001;
        mem[452] = 12'b000100100001;
        mem[453] = 12'b000100100010;
        mem[454] = 12'b000100100011;
        mem[455] = 12'b000100100011;
        mem[456] = 12'b000100100100;
        mem[457] = 12'b000100100100;
        mem[458] = 12'b000100100101;
        mem[459] = 12'b000100100110;
        mem[460] = 12'b000100100110;
        mem[461] = 12'b000100100111;
        mem[462] = 12'b000100101000;
        mem[463] = 12'b000100101000;
        mem[464] = 12'b000100101001;
        mem[465] = 12'b000100101010;
        mem[466] = 12'b000100101010;
        mem[467] = 12'b000100101011;
        mem[468] = 12'b000100101011;
        mem[469] = 12'b000100101100;
        mem[470] = 12'b000100101101;
        mem[471] = 12'b000100101101;
        mem[472] = 12'b000100101110;
        mem[473] = 12'b000100101111;
        mem[474] = 12'b000100101111;
        mem[475] = 12'b000100110000;
        mem[476] = 12'b000100110000;
        mem[477] = 12'b000100110001;
        mem[478] = 12'b000100110010;
        mem[479] = 12'b000100110010;
        mem[480] = 12'b000100110011;
        mem[481] = 12'b000100110100;
        mem[482] = 12'b000100110100;
        mem[483] = 12'b000100110101;
        mem[484] = 12'b000100110110;
        mem[485] = 12'b000100110110;
        mem[486] = 12'b000100110111;
        mem[487] = 12'b000100110111;
        mem[488] = 12'b000100111000;
        mem[489] = 12'b000100111001;
        mem[490] = 12'b000100111001;
        mem[491] = 12'b000100111010;
        mem[492] = 12'b000100111011;
        mem[493] = 12'b000100111011;
        mem[494] = 12'b000100111100;
        mem[495] = 12'b000100111101;
        mem[496] = 12'b000100111101;
        mem[497] = 12'b000100111110;
        mem[498] = 12'b000100111110;
        mem[499] = 12'b000100111111;
        mem[500] = 12'b000101000000;
        mem[501] = 12'b000101000000;
        mem[502] = 12'b000101000001;
        mem[503] = 12'b000101000010;
        mem[504] = 12'b000101000010;
        mem[505] = 12'b000101000011;
        mem[506] = 12'b000101000100;
        mem[507] = 12'b000101000100;
        mem[508] = 12'b000101000101;
        mem[509] = 12'b000101000101;
        mem[510] = 12'b000101000110;
        mem[511] = 12'b000101000111;
        mem[512] = 12'b000101000111;
        mem[513] = 12'b000101001000;
        mem[514] = 12'b000101001001;
        mem[515] = 12'b000101001001;
        mem[516] = 12'b000101001010;
        mem[517] = 12'b000101001011;
        mem[518] = 12'b000101001011;
        mem[519] = 12'b000101001100;
        mem[520] = 12'b000101001100;
        mem[521] = 12'b000101001101;
        mem[522] = 12'b000101001110;
        mem[523] = 12'b000101001110;
        mem[524] = 12'b000101001111;
        mem[525] = 12'b000101010000;
        mem[526] = 12'b000101010000;
        mem[527] = 12'b000101010001;
        mem[528] = 12'b000101010010;
        mem[529] = 12'b000101010010;
        mem[530] = 12'b000101010011;
        mem[531] = 12'b000101010011;
        mem[532] = 12'b000101010100;
        mem[533] = 12'b000101010101;
        mem[534] = 12'b000101010101;
        mem[535] = 12'b000101010110;
        mem[536] = 12'b000101010111;
        mem[537] = 12'b000101010111;
        mem[538] = 12'b000101011000;
        mem[539] = 12'b000101011001;
        mem[540] = 12'b000101011001;
        mem[541] = 12'b000101011010;
        mem[542] = 12'b000101011010;
        mem[543] = 12'b000101011011;
        mem[544] = 12'b000101011100;
        mem[545] = 12'b000101011100;
        mem[546] = 12'b000101011101;
        mem[547] = 12'b000101011110;
        mem[548] = 12'b000101011110;
        mem[549] = 12'b000101011111;
        mem[550] = 12'b000101011111;
        mem[551] = 12'b000101100000;
        mem[552] = 12'b000101100001;
        mem[553] = 12'b000101100001;
        mem[554] = 12'b000101100010;
        mem[555] = 12'b000101100011;
        mem[556] = 12'b000101100011;
        mem[557] = 12'b000101100100;
        mem[558] = 12'b000101100101;
        mem[559] = 12'b000101100101;
        mem[560] = 12'b000101100110;
        mem[561] = 12'b000101100110;
        mem[562] = 12'b000101100111;
        mem[563] = 12'b000101101000;
        mem[564] = 12'b000101101000;
        mem[565] = 12'b000101101001;
        mem[566] = 12'b000101101010;
        mem[567] = 12'b000101101010;
        mem[568] = 12'b000101101011;
        mem[569] = 12'b000101101100;
        mem[570] = 12'b000101101100;
        mem[571] = 12'b000101101101;
        mem[572] = 12'b000101101101;
        mem[573] = 12'b000101101110;
        mem[574] = 12'b000101101111;
        mem[575] = 12'b000101101111;
        mem[576] = 12'b000101110000;
        mem[577] = 12'b000101110001;
        mem[578] = 12'b000101110001;
        mem[579] = 12'b000101110010;
        mem[580] = 12'b000101110010;
        mem[581] = 12'b000101110011;
        mem[582] = 12'b000101110100;
        mem[583] = 12'b000101110100;
        mem[584] = 12'b000101110101;
        mem[585] = 12'b000101110110;
        mem[586] = 12'b000101110110;
        mem[587] = 12'b000101110111;
        mem[588] = 12'b000101111000;
        mem[589] = 12'b000101111000;
        mem[590] = 12'b000101111001;
        mem[591] = 12'b000101111001;
        mem[592] = 12'b000101111010;
        mem[593] = 12'b000101111011;
        mem[594] = 12'b000101111011;
        mem[595] = 12'b000101111100;
        mem[596] = 12'b000101111101;
        mem[597] = 12'b000101111101;
        mem[598] = 12'b000101111110;
        mem[599] = 12'b000101111110;
        mem[600] = 12'b000101111111;
        mem[601] = 12'b000110000000;
        mem[602] = 12'b000110000000;
        mem[603] = 12'b000110000001;
        mem[604] = 12'b000110000010;
        mem[605] = 12'b000110000010;
        mem[606] = 12'b000110000011;
        mem[607] = 12'b000110000100;
        mem[608] = 12'b000110000100;
        mem[609] = 12'b000110000101;
        mem[610] = 12'b000110000101;
        mem[611] = 12'b000110000110;
        mem[612] = 12'b000110000111;
        mem[613] = 12'b000110000111;
        mem[614] = 12'b000110001000;
        mem[615] = 12'b000110001001;
        mem[616] = 12'b000110001001;
        mem[617] = 12'b000110001010;
        mem[618] = 12'b000110001010;
        mem[619] = 12'b000110001011;
        mem[620] = 12'b000110001100;
        mem[621] = 12'b000110001100;
        mem[622] = 12'b000110001101;
        mem[623] = 12'b000110001110;
        mem[624] = 12'b000110001110;
        mem[625] = 12'b000110001111;
        mem[626] = 12'b000110010000;
        mem[627] = 12'b000110010000;
        mem[628] = 12'b000110010001;
        mem[629] = 12'b000110010001;
        mem[630] = 12'b000110010010;
        mem[631] = 12'b000110010011;
        mem[632] = 12'b000110010011;
        mem[633] = 12'b000110010100;
        mem[634] = 12'b000110010101;
        mem[635] = 12'b000110010101;
        mem[636] = 12'b000110010110;
        mem[637] = 12'b000110010110;
        mem[638] = 12'b000110010111;
        mem[639] = 12'b000110011000;
        mem[640] = 12'b000110011000;
        mem[641] = 12'b000110011001;
        mem[642] = 12'b000110011010;
        mem[643] = 12'b000110011010;
        mem[644] = 12'b000110011011;
        mem[645] = 12'b000110011011;
        mem[646] = 12'b000110011100;
        mem[647] = 12'b000110011101;
        mem[648] = 12'b000110011101;
        mem[649] = 12'b000110011110;
        mem[650] = 12'b000110011111;
        mem[651] = 12'b000110011111;
        mem[652] = 12'b000110100000;
        mem[653] = 12'b000110100001;
        mem[654] = 12'b000110100001;
        mem[655] = 12'b000110100010;
        mem[656] = 12'b000110100010;
        mem[657] = 12'b000110100011;
        mem[658] = 12'b000110100100;
        mem[659] = 12'b000110100100;
        mem[660] = 12'b000110100101;
        mem[661] = 12'b000110100110;
        mem[662] = 12'b000110100110;
        mem[663] = 12'b000110100111;
        mem[664] = 12'b000110100111;
        mem[665] = 12'b000110101000;
        mem[666] = 12'b000110101001;
        mem[667] = 12'b000110101001;
        mem[668] = 12'b000110101010;
        mem[669] = 12'b000110101011;
        mem[670] = 12'b000110101011;
        mem[671] = 12'b000110101100;
        mem[672] = 12'b000110101100;
        mem[673] = 12'b000110101101;
        mem[674] = 12'b000110101110;
        mem[675] = 12'b000110101110;
        mem[676] = 12'b000110101111;
        mem[677] = 12'b000110110000;
        mem[678] = 12'b000110110000;
        mem[679] = 12'b000110110001;
        mem[680] = 12'b000110110010;
        mem[681] = 12'b000110110010;
        mem[682] = 12'b000110110011;
        mem[683] = 12'b000110110011;
        mem[684] = 12'b000110110100;
        mem[685] = 12'b000110110101;
        mem[686] = 12'b000110110101;
        mem[687] = 12'b000110110110;
        mem[688] = 12'b000110110111;
        mem[689] = 12'b000110110111;
        mem[690] = 12'b000110111000;
        mem[691] = 12'b000110111000;
        mem[692] = 12'b000110111001;
        mem[693] = 12'b000110111010;
        mem[694] = 12'b000110111010;
        mem[695] = 12'b000110111011;
        mem[696] = 12'b000110111100;
        mem[697] = 12'b000110111100;
        mem[698] = 12'b000110111101;
        mem[699] = 12'b000110111101;
        mem[700] = 12'b000110111110;
        mem[701] = 12'b000110111111;
        mem[702] = 12'b000110111111;
        mem[703] = 12'b000111000000;
        mem[704] = 12'b000111000001;
        mem[705] = 12'b000111000001;
        mem[706] = 12'b000111000010;
        mem[707] = 12'b000111000010;
        mem[708] = 12'b000111000011;
        mem[709] = 12'b000111000100;
        mem[710] = 12'b000111000100;
        mem[711] = 12'b000111000101;
        mem[712] = 12'b000111000110;
        mem[713] = 12'b000111000110;
        mem[714] = 12'b000111000111;
        mem[715] = 12'b000111000111;
        mem[716] = 12'b000111001000;
        mem[717] = 12'b000111001001;
        mem[718] = 12'b000111001001;
        mem[719] = 12'b000111001010;
        mem[720] = 12'b000111001011;
        mem[721] = 12'b000111001011;
        mem[722] = 12'b000111001100;
        mem[723] = 12'b000111001101;
        mem[724] = 12'b000111001101;
        mem[725] = 12'b000111001110;
        mem[726] = 12'b000111001110;
        mem[727] = 12'b000111001111;
        mem[728] = 12'b000111010000;
        mem[729] = 12'b000111010000;
        mem[730] = 12'b000111010001;
        mem[731] = 12'b000111010010;
        mem[732] = 12'b000111010010;
        mem[733] = 12'b000111010011;
        mem[734] = 12'b000111010011;
        mem[735] = 12'b000111010100;
        mem[736] = 12'b000111010101;
        mem[737] = 12'b000111010101;
        mem[738] = 12'b000111010110;
        mem[739] = 12'b000111010111;
        mem[740] = 12'b000111010111;
        mem[741] = 12'b000111011000;
        mem[742] = 12'b000111011000;
        mem[743] = 12'b000111011001;
        mem[744] = 12'b000111011010;
        mem[745] = 12'b000111011010;
        mem[746] = 12'b000111011011;
        mem[747] = 12'b000111011100;
        mem[748] = 12'b000111011100;
        mem[749] = 12'b000111011101;
        mem[750] = 12'b000111011101;
        mem[751] = 12'b000111011110;
        mem[752] = 12'b000111011111;
        mem[753] = 12'b000111011111;
        mem[754] = 12'b000111100000;
        mem[755] = 12'b000111100001;
        mem[756] = 12'b000111100001;
        mem[757] = 12'b000111100010;
        mem[758] = 12'b000111100010;
        mem[759] = 12'b000111100011;
        mem[760] = 12'b000111100100;
        mem[761] = 12'b000111100100;
        mem[762] = 12'b000111100101;
        mem[763] = 12'b000111100110;
        mem[764] = 12'b000111100110;
        mem[765] = 12'b000111100111;
        mem[766] = 12'b000111100111;
        mem[767] = 12'b000111101000;
        mem[768] = 12'b000111101001;
        mem[769] = 12'b000111101001;
        mem[770] = 12'b000111101010;
        mem[771] = 12'b000111101011;
        mem[772] = 12'b000111101011;
        mem[773] = 12'b000111101100;
        mem[774] = 12'b000111101100;
        mem[775] = 12'b000111101101;
        mem[776] = 12'b000111101110;
        mem[777] = 12'b000111101110;
        mem[778] = 12'b000111101111;
        mem[779] = 12'b000111110000;
        mem[780] = 12'b000111110000;
        mem[781] = 12'b000111110001;
        mem[782] = 12'b000111110001;
        mem[783] = 12'b000111110010;
        mem[784] = 12'b000111110011;
        mem[785] = 12'b000111110011;
        mem[786] = 12'b000111110100;
        mem[787] = 12'b000111110101;
        mem[788] = 12'b000111110101;
        mem[789] = 12'b000111110110;
        mem[790] = 12'b000111110110;
        mem[791] = 12'b000111110111;
        mem[792] = 12'b000111111000;
        mem[793] = 12'b000111111000;
        mem[794] = 12'b000111111001;
        mem[795] = 12'b000111111010;
        mem[796] = 12'b000111111010;
        mem[797] = 12'b000111111011;
        mem[798] = 12'b000111111011;
        mem[799] = 12'b000111111100;
        mem[800] = 12'b000111111101;
        mem[801] = 12'b000111111101;
        mem[802] = 12'b000111111110;
        mem[803] = 12'b000111111110;
        mem[804] = 12'b000111111111;
        mem[805] = 12'b001000000000;
        mem[806] = 12'b001000000000;
        mem[807] = 12'b001000000001;
        mem[808] = 12'b001000000010;
        mem[809] = 12'b001000000010;
        mem[810] = 12'b001000000011;
        mem[811] = 12'b001000000011;
        mem[812] = 12'b001000000100;
        mem[813] = 12'b001000000101;
        mem[814] = 12'b001000000101;
        mem[815] = 12'b001000000110;
        mem[816] = 12'b001000000111;
        mem[817] = 12'b001000000111;
        mem[818] = 12'b001000001000;
        mem[819] = 12'b001000001000;
        mem[820] = 12'b001000001001;
        mem[821] = 12'b001000001010;
        mem[822] = 12'b001000001010;
        mem[823] = 12'b001000001011;
        mem[824] = 12'b001000001100;
        mem[825] = 12'b001000001100;
        mem[826] = 12'b001000001101;
        mem[827] = 12'b001000001101;
        mem[828] = 12'b001000001110;
        mem[829] = 12'b001000001111;
        mem[830] = 12'b001000001111;
        mem[831] = 12'b001000010000;
        mem[832] = 12'b001000010001;
        mem[833] = 12'b001000010001;
        mem[834] = 12'b001000010010;
        mem[835] = 12'b001000010010;
        mem[836] = 12'b001000010011;
        mem[837] = 12'b001000010100;
        mem[838] = 12'b001000010100;
        mem[839] = 12'b001000010101;
        mem[840] = 12'b001000010101;
        mem[841] = 12'b001000010110;
        mem[842] = 12'b001000010111;
        mem[843] = 12'b001000010111;
        mem[844] = 12'b001000011000;
        mem[845] = 12'b001000011001;
        mem[846] = 12'b001000011001;
        mem[847] = 12'b001000011010;
        mem[848] = 12'b001000011010;
        mem[849] = 12'b001000011011;
        mem[850] = 12'b001000011100;
        mem[851] = 12'b001000011100;
        mem[852] = 12'b001000011101;
        mem[853] = 12'b001000011110;
        mem[854] = 12'b001000011110;
        mem[855] = 12'b001000011111;
        mem[856] = 12'b001000011111;
        mem[857] = 12'b001000100000;
        mem[858] = 12'b001000100001;
        mem[859] = 12'b001000100001;
        mem[860] = 12'b001000100010;
        mem[861] = 12'b001000100011;
        mem[862] = 12'b001000100011;
        mem[863] = 12'b001000100100;
        mem[864] = 12'b001000100100;
        mem[865] = 12'b001000100101;
        mem[866] = 12'b001000100110;
        mem[867] = 12'b001000100110;
        mem[868] = 12'b001000100111;
        mem[869] = 12'b001000100111;
        mem[870] = 12'b001000101000;
        mem[871] = 12'b001000101001;
        mem[872] = 12'b001000101001;
        mem[873] = 12'b001000101010;
        mem[874] = 12'b001000101011;
        mem[875] = 12'b001000101011;
        mem[876] = 12'b001000101100;
        mem[877] = 12'b001000101100;
        mem[878] = 12'b001000101101;
        mem[879] = 12'b001000101110;
        mem[880] = 12'b001000101110;
        mem[881] = 12'b001000101111;
        mem[882] = 12'b001000110000;
        mem[883] = 12'b001000110000;
        mem[884] = 12'b001000110001;
        mem[885] = 12'b001000110001;
        mem[886] = 12'b001000110010;
        mem[887] = 12'b001000110011;
        mem[888] = 12'b001000110011;
        mem[889] = 12'b001000110100;
        mem[890] = 12'b001000110100;
        mem[891] = 12'b001000110101;
        mem[892] = 12'b001000110110;
        mem[893] = 12'b001000110110;
        mem[894] = 12'b001000110111;
        mem[895] = 12'b001000111000;
        mem[896] = 12'b001000111000;
        mem[897] = 12'b001000111001;
        mem[898] = 12'b001000111001;
        mem[899] = 12'b001000111010;
        mem[900] = 12'b001000111011;
        mem[901] = 12'b001000111011;
        mem[902] = 12'b001000111100;
        mem[903] = 12'b001000111101;
        mem[904] = 12'b001000111101;
        mem[905] = 12'b001000111110;
        mem[906] = 12'b001000111110;
        mem[907] = 12'b001000111111;
        mem[908] = 12'b001001000000;
        mem[909] = 12'b001001000000;
        mem[910] = 12'b001001000001;
        mem[911] = 12'b001001000001;
        mem[912] = 12'b001001000010;
        mem[913] = 12'b001001000011;
        mem[914] = 12'b001001000011;
        mem[915] = 12'b001001000100;
        mem[916] = 12'b001001000101;
        mem[917] = 12'b001001000101;
        mem[918] = 12'b001001000110;
        mem[919] = 12'b001001000110;
        mem[920] = 12'b001001000111;
        mem[921] = 12'b001001001000;
        mem[922] = 12'b001001001000;
        mem[923] = 12'b001001001001;
        mem[924] = 12'b001001001001;
        mem[925] = 12'b001001001010;
        mem[926] = 12'b001001001011;
        mem[927] = 12'b001001001011;
        mem[928] = 12'b001001001100;
        mem[929] = 12'b001001001101;
        mem[930] = 12'b001001001101;
        mem[931] = 12'b001001001110;
        mem[932] = 12'b001001001110;
        mem[933] = 12'b001001001111;
        mem[934] = 12'b001001010000;
        mem[935] = 12'b001001010000;
        mem[936] = 12'b001001010001;
        mem[937] = 12'b001001010001;
        mem[938] = 12'b001001010010;
        mem[939] = 12'b001001010011;
        mem[940] = 12'b001001010011;
        mem[941] = 12'b001001010100;
        mem[942] = 12'b001001010101;
        mem[943] = 12'b001001010101;
        mem[944] = 12'b001001010110;
        mem[945] = 12'b001001010110;
        mem[946] = 12'b001001010111;
        mem[947] = 12'b001001011000;
        mem[948] = 12'b001001011000;
        mem[949] = 12'b001001011001;
        mem[950] = 12'b001001011001;
        mem[951] = 12'b001001011010;
        mem[952] = 12'b001001011011;
        mem[953] = 12'b001001011011;
        mem[954] = 12'b001001011100;
        mem[955] = 12'b001001011101;
        mem[956] = 12'b001001011101;
        mem[957] = 12'b001001011110;
        mem[958] = 12'b001001011110;
        mem[959] = 12'b001001011111;
        mem[960] = 12'b001001100000;
        mem[961] = 12'b001001100000;
        mem[962] = 12'b001001100001;
        mem[963] = 12'b001001100001;
        mem[964] = 12'b001001100010;
        mem[965] = 12'b001001100011;
        mem[966] = 12'b001001100011;
        mem[967] = 12'b001001100100;
        mem[968] = 12'b001001100101;
        mem[969] = 12'b001001100101;
        mem[970] = 12'b001001100110;
        mem[971] = 12'b001001100110;
        mem[972] = 12'b001001100111;
        mem[973] = 12'b001001101000;
        mem[974] = 12'b001001101000;
        mem[975] = 12'b001001101001;
        mem[976] = 12'b001001101001;
        mem[977] = 12'b001001101010;
        mem[978] = 12'b001001101011;
        mem[979] = 12'b001001101011;
        mem[980] = 12'b001001101100;
        mem[981] = 12'b001001101100;
        mem[982] = 12'b001001101101;
        mem[983] = 12'b001001101110;
        mem[984] = 12'b001001101110;
        mem[985] = 12'b001001101111;
        mem[986] = 12'b001001110000;
        mem[987] = 12'b001001110000;
        mem[988] = 12'b001001110001;
        mem[989] = 12'b001001110001;
        mem[990] = 12'b001001110010;
        mem[991] = 12'b001001110011;
        mem[992] = 12'b001001110011;
        mem[993] = 12'b001001110100;
        mem[994] = 12'b001001110100;
        mem[995] = 12'b001001110101;
        mem[996] = 12'b001001110110;
        mem[997] = 12'b001001110110;
        mem[998] = 12'b001001110111;
        mem[999] = 12'b001001111000;
        mem[1000] = 12'b001001111000;
        mem[1001] = 12'b001001111001;
        mem[1002] = 12'b001001111001;
        mem[1003] = 12'b001001111010;
        mem[1004] = 12'b001001111011;
        mem[1005] = 12'b001001111011;
        mem[1006] = 12'b001001111100;
        mem[1007] = 12'b001001111100;
        mem[1008] = 12'b001001111101;
        mem[1009] = 12'b001001111110;
        mem[1010] = 12'b001001111110;
        mem[1011] = 12'b001001111111;
        mem[1012] = 12'b001001111111;
        mem[1013] = 12'b001010000000;
        mem[1014] = 12'b001010000001;
        mem[1015] = 12'b001010000001;
        mem[1016] = 12'b001010000010;
        mem[1017] = 12'b001010000011;
        mem[1018] = 12'b001010000011;
        mem[1019] = 12'b001010000100;
        mem[1020] = 12'b001010000100;
        mem[1021] = 12'b001010000101;
        mem[1022] = 12'b001010000110;
        mem[1023] = 12'b001010000110;
        mem[1024] = 12'b001010000111;
        mem[1025] = 12'b001010000111;
        mem[1026] = 12'b001010001000;
        mem[1027] = 12'b001010001001;
        mem[1028] = 12'b001010001001;
        mem[1029] = 12'b001010001010;
        mem[1030] = 12'b001010001010;
        mem[1031] = 12'b001010001011;
        mem[1032] = 12'b001010001100;
        mem[1033] = 12'b001010001100;
        mem[1034] = 12'b001010001101;
        mem[1035] = 12'b001010001101;
        mem[1036] = 12'b001010001110;
        mem[1037] = 12'b001010001111;
        mem[1038] = 12'b001010001111;
        mem[1039] = 12'b001010010000;
        mem[1040] = 12'b001010010001;
        mem[1041] = 12'b001010010001;
        mem[1042] = 12'b001010010010;
        mem[1043] = 12'b001010010010;
        mem[1044] = 12'b001010010011;
        mem[1045] = 12'b001010010100;
        mem[1046] = 12'b001010010100;
        mem[1047] = 12'b001010010101;
        mem[1048] = 12'b001010010101;
        mem[1049] = 12'b001010010110;
        mem[1050] = 12'b001010010111;
        mem[1051] = 12'b001010010111;
        mem[1052] = 12'b001010011000;
        mem[1053] = 12'b001010011000;
        mem[1054] = 12'b001010011001;
        mem[1055] = 12'b001010011010;
        mem[1056] = 12'b001010011010;
        mem[1057] = 12'b001010011011;
        mem[1058] = 12'b001010011011;
        mem[1059] = 12'b001010011100;
        mem[1060] = 12'b001010011101;
        mem[1061] = 12'b001010011101;
        mem[1062] = 12'b001010011110;
        mem[1063] = 12'b001010011111;
        mem[1064] = 12'b001010011111;
        mem[1065] = 12'b001010100000;
        mem[1066] = 12'b001010100000;
        mem[1067] = 12'b001010100001;
        mem[1068] = 12'b001010100010;
        mem[1069] = 12'b001010100010;
        mem[1070] = 12'b001010100011;
        mem[1071] = 12'b001010100011;
        mem[1072] = 12'b001010100100;
        mem[1073] = 12'b001010100101;
        mem[1074] = 12'b001010100101;
        mem[1075] = 12'b001010100110;
        mem[1076] = 12'b001010100110;
        mem[1077] = 12'b001010100111;
        mem[1078] = 12'b001010101000;
        mem[1079] = 12'b001010101000;
        mem[1080] = 12'b001010101001;
        mem[1081] = 12'b001010101001;
        mem[1082] = 12'b001010101010;
        mem[1083] = 12'b001010101011;
        mem[1084] = 12'b001010101011;
        mem[1085] = 12'b001010101100;
        mem[1086] = 12'b001010101100;
        mem[1087] = 12'b001010101101;
        mem[1088] = 12'b001010101110;
        mem[1089] = 12'b001010101110;
        mem[1090] = 12'b001010101111;
        mem[1091] = 12'b001010110000;
        mem[1092] = 12'b001010110000;
        mem[1093] = 12'b001010110001;
        mem[1094] = 12'b001010110001;
        mem[1095] = 12'b001010110010;
        mem[1096] = 12'b001010110011;
        mem[1097] = 12'b001010110011;
        mem[1098] = 12'b001010110100;
        mem[1099] = 12'b001010110100;
        mem[1100] = 12'b001010110101;
        mem[1101] = 12'b001010110110;
        mem[1102] = 12'b001010110110;
        mem[1103] = 12'b001010110111;
        mem[1104] = 12'b001010110111;
        mem[1105] = 12'b001010111000;
        mem[1106] = 12'b001010111001;
        mem[1107] = 12'b001010111001;
        mem[1108] = 12'b001010111010;
        mem[1109] = 12'b001010111010;
        mem[1110] = 12'b001010111011;
        mem[1111] = 12'b001010111100;
        mem[1112] = 12'b001010111100;
        mem[1113] = 12'b001010111101;
        mem[1114] = 12'b001010111101;
        mem[1115] = 12'b001010111110;
        mem[1116] = 12'b001010111111;
        mem[1117] = 12'b001010111111;
        mem[1118] = 12'b001011000000;
        mem[1119] = 12'b001011000000;
        mem[1120] = 12'b001011000001;
        mem[1121] = 12'b001011000010;
        mem[1122] = 12'b001011000010;
        mem[1123] = 12'b001011000011;
        mem[1124] = 12'b001011000011;
        mem[1125] = 12'b001011000100;
        mem[1126] = 12'b001011000101;
        mem[1127] = 12'b001011000101;
        mem[1128] = 12'b001011000110;
        mem[1129] = 12'b001011000110;
        mem[1130] = 12'b001011000111;
        mem[1131] = 12'b001011001000;
        mem[1132] = 12'b001011001000;
        mem[1133] = 12'b001011001001;
        mem[1134] = 12'b001011001001;
        mem[1135] = 12'b001011001010;
        mem[1136] = 12'b001011001011;
        mem[1137] = 12'b001011001011;
        mem[1138] = 12'b001011001100;
        mem[1139] = 12'b001011001101;
        mem[1140] = 12'b001011001101;
        mem[1141] = 12'b001011001110;
        mem[1142] = 12'b001011001110;
        mem[1143] = 12'b001011001111;
        mem[1144] = 12'b001011010000;
        mem[1145] = 12'b001011010000;
        mem[1146] = 12'b001011010001;
        mem[1147] = 12'b001011010001;
        mem[1148] = 12'b001011010010;
        mem[1149] = 12'b001011010011;
        mem[1150] = 12'b001011010011;
        mem[1151] = 12'b001011010100;
        mem[1152] = 12'b001011010100;
        mem[1153] = 12'b001011010101;
        mem[1154] = 12'b001011010110;
        mem[1155] = 12'b001011010110;
        mem[1156] = 12'b001011010111;
        mem[1157] = 12'b001011010111;
        mem[1158] = 12'b001011011000;
        mem[1159] = 12'b001011011001;
        mem[1160] = 12'b001011011001;
        mem[1161] = 12'b001011011010;
        mem[1162] = 12'b001011011010;
        mem[1163] = 12'b001011011011;
        mem[1164] = 12'b001011011100;
        mem[1165] = 12'b001011011100;
        mem[1166] = 12'b001011011101;
        mem[1167] = 12'b001011011101;
        mem[1168] = 12'b001011011110;
        mem[1169] = 12'b001011011111;
        mem[1170] = 12'b001011011111;
        mem[1171] = 12'b001011100000;
        mem[1172] = 12'b001011100000;
        mem[1173] = 12'b001011100001;
        mem[1174] = 12'b001011100010;
        mem[1175] = 12'b001011100010;
        mem[1176] = 12'b001011100011;
        mem[1177] = 12'b001011100011;
        mem[1178] = 12'b001011100100;
        mem[1179] = 12'b001011100101;
        mem[1180] = 12'b001011100101;
        mem[1181] = 12'b001011100110;
        mem[1182] = 12'b001011100110;
        mem[1183] = 12'b001011100111;
        mem[1184] = 12'b001011101000;
        mem[1185] = 12'b001011101000;
        mem[1186] = 12'b001011101001;
        mem[1187] = 12'b001011101001;
        mem[1188] = 12'b001011101010;
        mem[1189] = 12'b001011101011;
        mem[1190] = 12'b001011101011;
        mem[1191] = 12'b001011101100;
        mem[1192] = 12'b001011101100;
        mem[1193] = 12'b001011101101;
        mem[1194] = 12'b001011101110;
        mem[1195] = 12'b001011101110;
        mem[1196] = 12'b001011101111;
        mem[1197] = 12'b001011101111;
        mem[1198] = 12'b001011110000;
        mem[1199] = 12'b001011110001;
        mem[1200] = 12'b001011110001;
        mem[1201] = 12'b001011110010;
        mem[1202] = 12'b001011110010;
        mem[1203] = 12'b001011110011;
        mem[1204] = 12'b001011110100;
        mem[1205] = 12'b001011110100;
        mem[1206] = 12'b001011110101;
        mem[1207] = 12'b001011110101;
        mem[1208] = 12'b001011110110;
        mem[1209] = 12'b001011110111;
        mem[1210] = 12'b001011110111;
        mem[1211] = 12'b001011111000;
        mem[1212] = 12'b001011111000;
        mem[1213] = 12'b001011111001;
        mem[1214] = 12'b001011111001;
        mem[1215] = 12'b001011111010;
        mem[1216] = 12'b001011111011;
        mem[1217] = 12'b001011111011;
        mem[1218] = 12'b001011111100;
        mem[1219] = 12'b001011111100;
        mem[1220] = 12'b001011111101;
        mem[1221] = 12'b001011111110;
        mem[1222] = 12'b001011111110;
        mem[1223] = 12'b001011111111;
        mem[1224] = 12'b001011111111;
        mem[1225] = 12'b001100000000;
        mem[1226] = 12'b001100000001;
        mem[1227] = 12'b001100000001;
        mem[1228] = 12'b001100000010;
        mem[1229] = 12'b001100000010;
        mem[1230] = 12'b001100000011;
        mem[1231] = 12'b001100000100;
        mem[1232] = 12'b001100000100;
        mem[1233] = 12'b001100000101;
        mem[1234] = 12'b001100000101;
        mem[1235] = 12'b001100000110;
        mem[1236] = 12'b001100000111;
        mem[1237] = 12'b001100000111;
        mem[1238] = 12'b001100001000;
        mem[1239] = 12'b001100001000;
        mem[1240] = 12'b001100001001;
        mem[1241] = 12'b001100001010;
        mem[1242] = 12'b001100001010;
        mem[1243] = 12'b001100001011;
        mem[1244] = 12'b001100001011;
        mem[1245] = 12'b001100001100;
        mem[1246] = 12'b001100001101;
        mem[1247] = 12'b001100001101;
        mem[1248] = 12'b001100001110;
        mem[1249] = 12'b001100001110;
        mem[1250] = 12'b001100001111;
        mem[1251] = 12'b001100010000;
        mem[1252] = 12'b001100010000;
        mem[1253] = 12'b001100010001;
        mem[1254] = 12'b001100010001;
        mem[1255] = 12'b001100010010;
        mem[1256] = 12'b001100010010;
        mem[1257] = 12'b001100010011;
        mem[1258] = 12'b001100010100;
        mem[1259] = 12'b001100010100;
        mem[1260] = 12'b001100010101;
        mem[1261] = 12'b001100010101;
        mem[1262] = 12'b001100010110;
        mem[1263] = 12'b001100010111;
        mem[1264] = 12'b001100010111;
        mem[1265] = 12'b001100011000;
        mem[1266] = 12'b001100011000;
        mem[1267] = 12'b001100011001;
        mem[1268] = 12'b001100011010;
        mem[1269] = 12'b001100011010;
        mem[1270] = 12'b001100011011;
        mem[1271] = 12'b001100011011;
        mem[1272] = 12'b001100011100;
        mem[1273] = 12'b001100011101;
        mem[1274] = 12'b001100011101;
        mem[1275] = 12'b001100011110;
        mem[1276] = 12'b001100011110;
        mem[1277] = 12'b001100011111;
        mem[1278] = 12'b001100100000;
        mem[1279] = 12'b001100100000;
        mem[1280] = 12'b001100100001;
        mem[1281] = 12'b001100100001;
        mem[1282] = 12'b001100100010;
        mem[1283] = 12'b001100100010;
        mem[1284] = 12'b001100100011;
        mem[1285] = 12'b001100100100;
        mem[1286] = 12'b001100100100;
        mem[1287] = 12'b001100100101;
        mem[1288] = 12'b001100100101;
        mem[1289] = 12'b001100100110;
        mem[1290] = 12'b001100100111;
        mem[1291] = 12'b001100100111;
        mem[1292] = 12'b001100101000;
        mem[1293] = 12'b001100101000;
        mem[1294] = 12'b001100101001;
        mem[1295] = 12'b001100101010;
        mem[1296] = 12'b001100101010;
        mem[1297] = 12'b001100101011;
        mem[1298] = 12'b001100101011;
        mem[1299] = 12'b001100101100;
        mem[1300] = 12'b001100101101;
        mem[1301] = 12'b001100101101;
        mem[1302] = 12'b001100101110;
        mem[1303] = 12'b001100101110;
        mem[1304] = 12'b001100101111;
        mem[1305] = 12'b001100101111;
        mem[1306] = 12'b001100110000;
        mem[1307] = 12'b001100110001;
        mem[1308] = 12'b001100110001;
        mem[1309] = 12'b001100110010;
        mem[1310] = 12'b001100110010;
        mem[1311] = 12'b001100110011;
        mem[1312] = 12'b001100110100;
        mem[1313] = 12'b001100110100;
        mem[1314] = 12'b001100110101;
        mem[1315] = 12'b001100110101;
        mem[1316] = 12'b001100110110;
        mem[1317] = 12'b001100110111;
        mem[1318] = 12'b001100110111;
        mem[1319] = 12'b001100111000;
        mem[1320] = 12'b001100111000;
        mem[1321] = 12'b001100111001;
        mem[1322] = 12'b001100111010;
        mem[1323] = 12'b001100111010;
        mem[1324] = 12'b001100111011;
        mem[1325] = 12'b001100111011;
        mem[1326] = 12'b001100111100;
        mem[1327] = 12'b001100111100;
        mem[1328] = 12'b001100111101;
        mem[1329] = 12'b001100111110;
        mem[1330] = 12'b001100111110;
        mem[1331] = 12'b001100111111;
        mem[1332] = 12'b001100111111;
        mem[1333] = 12'b001101000000;
        mem[1334] = 12'b001101000001;
        mem[1335] = 12'b001101000001;
        mem[1336] = 12'b001101000010;
        mem[1337] = 12'b001101000010;
        mem[1338] = 12'b001101000011;
        mem[1339] = 12'b001101000011;
        mem[1340] = 12'b001101000100;
        mem[1341] = 12'b001101000101;
        mem[1342] = 12'b001101000101;
        mem[1343] = 12'b001101000110;
        mem[1344] = 12'b001101000110;
        mem[1345] = 12'b001101000111;
        mem[1346] = 12'b001101001000;
        mem[1347] = 12'b001101001000;
        mem[1348] = 12'b001101001001;
        mem[1349] = 12'b001101001001;
        mem[1350] = 12'b001101001010;
        mem[1351] = 12'b001101001011;
        mem[1352] = 12'b001101001011;
        mem[1353] = 12'b001101001100;
        mem[1354] = 12'b001101001100;
        mem[1355] = 12'b001101001101;
        mem[1356] = 12'b001101001101;
        mem[1357] = 12'b001101001110;
        mem[1358] = 12'b001101001111;
        mem[1359] = 12'b001101001111;
        mem[1360] = 12'b001101010000;
        mem[1361] = 12'b001101010000;
        mem[1362] = 12'b001101010001;
        mem[1363] = 12'b001101010010;
        mem[1364] = 12'b001101010010;
        mem[1365] = 12'b001101010011;
        mem[1366] = 12'b001101010011;
        mem[1367] = 12'b001101010100;
        mem[1368] = 12'b001101010100;
        mem[1369] = 12'b001101010101;
        mem[1370] = 12'b001101010110;
        mem[1371] = 12'b001101010110;
        mem[1372] = 12'b001101010111;
        mem[1373] = 12'b001101010111;
        mem[1374] = 12'b001101011000;
        mem[1375] = 12'b001101011001;
        mem[1376] = 12'b001101011001;
        mem[1377] = 12'b001101011010;
        mem[1378] = 12'b001101011010;
        mem[1379] = 12'b001101011011;
        mem[1380] = 12'b001101011011;
        mem[1381] = 12'b001101011100;
        mem[1382] = 12'b001101011101;
        mem[1383] = 12'b001101011101;
        mem[1384] = 12'b001101011110;
        mem[1385] = 12'b001101011110;
        mem[1386] = 12'b001101011111;
        mem[1387] = 12'b001101100000;
        mem[1388] = 12'b001101100000;
        mem[1389] = 12'b001101100001;
        mem[1390] = 12'b001101100001;
        mem[1391] = 12'b001101100010;
        mem[1392] = 12'b001101100010;
        mem[1393] = 12'b001101100011;
        mem[1394] = 12'b001101100100;
        mem[1395] = 12'b001101100100;
        mem[1396] = 12'b001101100101;
        mem[1397] = 12'b001101100101;
        mem[1398] = 12'b001101100110;
        mem[1399] = 12'b001101100111;
        mem[1400] = 12'b001101100111;
        mem[1401] = 12'b001101101000;
        mem[1402] = 12'b001101101000;
        mem[1403] = 12'b001101101001;
        mem[1404] = 12'b001101101001;
        mem[1405] = 12'b001101101010;
        mem[1406] = 12'b001101101011;
        mem[1407] = 12'b001101101011;
        mem[1408] = 12'b001101101100;
        mem[1409] = 12'b001101101100;
        mem[1410] = 12'b001101101101;
        mem[1411] = 12'b001101101110;
        mem[1412] = 12'b001101101110;
        mem[1413] = 12'b001101101111;
        mem[1414] = 12'b001101101111;
        mem[1415] = 12'b001101110000;
        mem[1416] = 12'b001101110000;
        mem[1417] = 12'b001101110001;
        mem[1418] = 12'b001101110010;
        mem[1419] = 12'b001101110010;
        mem[1420] = 12'b001101110011;
        mem[1421] = 12'b001101110011;
        mem[1422] = 12'b001101110100;
        mem[1423] = 12'b001101110101;
        mem[1424] = 12'b001101110101;
        mem[1425] = 12'b001101110110;
        mem[1426] = 12'b001101110110;
        mem[1427] = 12'b001101110111;
        mem[1428] = 12'b001101110111;
        mem[1429] = 12'b001101111000;
        mem[1430] = 12'b001101111001;
        mem[1431] = 12'b001101111001;
        mem[1432] = 12'b001101111010;
        mem[1433] = 12'b001101111010;
        mem[1434] = 12'b001101111011;
        mem[1435] = 12'b001101111011;
        mem[1436] = 12'b001101111100;
        mem[1437] = 12'b001101111101;
        mem[1438] = 12'b001101111101;
        mem[1439] = 12'b001101111110;
        mem[1440] = 12'b001101111110;
        mem[1441] = 12'b001101111111;
        mem[1442] = 12'b001110000000;
        mem[1443] = 12'b001110000000;
        mem[1444] = 12'b001110000001;
        mem[1445] = 12'b001110000001;
        mem[1446] = 12'b001110000010;
        mem[1447] = 12'b001110000010;
        mem[1448] = 12'b001110000011;
        mem[1449] = 12'b001110000100;
        mem[1450] = 12'b001110000100;
        mem[1451] = 12'b001110000101;
        mem[1452] = 12'b001110000101;
        mem[1453] = 12'b001110000110;
        mem[1454] = 12'b001110000110;
        mem[1455] = 12'b001110000111;
        mem[1456] = 12'b001110001000;
        mem[1457] = 12'b001110001000;
        mem[1458] = 12'b001110001001;
        mem[1459] = 12'b001110001001;
        mem[1460] = 12'b001110001010;
        mem[1461] = 12'b001110001010;
        mem[1462] = 12'b001110001011;
        mem[1463] = 12'b001110001100;
        mem[1464] = 12'b001110001100;
        mem[1465] = 12'b001110001101;
        mem[1466] = 12'b001110001101;
        mem[1467] = 12'b001110001110;
        mem[1468] = 12'b001110001111;
        mem[1469] = 12'b001110001111;
        mem[1470] = 12'b001110010000;
        mem[1471] = 12'b001110010000;
        mem[1472] = 12'b001110010001;
        mem[1473] = 12'b001110010001;
        mem[1474] = 12'b001110010010;
        mem[1475] = 12'b001110010011;
        mem[1476] = 12'b001110010011;
        mem[1477] = 12'b001110010100;
        mem[1478] = 12'b001110010100;
        mem[1479] = 12'b001110010101;
        mem[1480] = 12'b001110010101;
        mem[1481] = 12'b001110010110;
        mem[1482] = 12'b001110010111;
        mem[1483] = 12'b001110010111;
        mem[1484] = 12'b001110011000;
        mem[1485] = 12'b001110011000;
        mem[1486] = 12'b001110011001;
        mem[1487] = 12'b001110011001;
        mem[1488] = 12'b001110011010;
        mem[1489] = 12'b001110011011;
        mem[1490] = 12'b001110011011;
        mem[1491] = 12'b001110011100;
        mem[1492] = 12'b001110011100;
        mem[1493] = 12'b001110011101;
        mem[1494] = 12'b001110011101;
        mem[1495] = 12'b001110011110;
        mem[1496] = 12'b001110011111;
        mem[1497] = 12'b001110011111;
        mem[1498] = 12'b001110100000;
        mem[1499] = 12'b001110100000;
        mem[1500] = 12'b001110100001;
        mem[1501] = 12'b001110100001;
        mem[1502] = 12'b001110100010;
        mem[1503] = 12'b001110100011;
        mem[1504] = 12'b001110100011;
        mem[1505] = 12'b001110100100;
        mem[1506] = 12'b001110100100;
        mem[1507] = 12'b001110100101;
        mem[1508] = 12'b001110100101;
        mem[1509] = 12'b001110100110;
        mem[1510] = 12'b001110100111;
        mem[1511] = 12'b001110100111;
        mem[1512] = 12'b001110101000;
        mem[1513] = 12'b001110101000;
        mem[1514] = 12'b001110101001;
        mem[1515] = 12'b001110101001;
        mem[1516] = 12'b001110101010;
        mem[1517] = 12'b001110101011;
        mem[1518] = 12'b001110101011;
        mem[1519] = 12'b001110101100;
        mem[1520] = 12'b001110101100;
        mem[1521] = 12'b001110101101;
        mem[1522] = 12'b001110101101;
        mem[1523] = 12'b001110101110;
        mem[1524] = 12'b001110101111;
        mem[1525] = 12'b001110101111;
        mem[1526] = 12'b001110110000;
        mem[1527] = 12'b001110110000;
        mem[1528] = 12'b001110110001;
        mem[1529] = 12'b001110110001;
        mem[1530] = 12'b001110110010;
        mem[1531] = 12'b001110110011;
        mem[1532] = 12'b001110110011;
        mem[1533] = 12'b001110110100;
        mem[1534] = 12'b001110110100;
        mem[1535] = 12'b001110110101;
        mem[1536] = 12'b001110110101;
        mem[1537] = 12'b001110110110;
        mem[1538] = 12'b001110110111;
        mem[1539] = 12'b001110110111;
        mem[1540] = 12'b001110111000;
        mem[1541] = 12'b001110111000;
        mem[1542] = 12'b001110111001;
        mem[1543] = 12'b001110111001;
        mem[1544] = 12'b001110111010;
        mem[1545] = 12'b001110111011;
        mem[1546] = 12'b001110111011;
        mem[1547] = 12'b001110111100;
        mem[1548] = 12'b001110111100;
        mem[1549] = 12'b001110111101;
        mem[1550] = 12'b001110111101;
        mem[1551] = 12'b001110111110;
        mem[1552] = 12'b001110111111;
        mem[1553] = 12'b001110111111;
        mem[1554] = 12'b001111000000;
        mem[1555] = 12'b001111000000;
        mem[1556] = 12'b001111000001;
        mem[1557] = 12'b001111000001;
        mem[1558] = 12'b001111000010;
        mem[1559] = 12'b001111000011;
        mem[1560] = 12'b001111000011;
        mem[1561] = 12'b001111000100;
        mem[1562] = 12'b001111000100;
        mem[1563] = 12'b001111000101;
        mem[1564] = 12'b001111000101;
        mem[1565] = 12'b001111000110;
        mem[1566] = 12'b001111000111;
        mem[1567] = 12'b001111000111;
        mem[1568] = 12'b001111001000;
        mem[1569] = 12'b001111001000;
        mem[1570] = 12'b001111001001;
        mem[1571] = 12'b001111001001;
        mem[1572] = 12'b001111001010;
        mem[1573] = 12'b001111001010;
        mem[1574] = 12'b001111001011;
        mem[1575] = 12'b001111001100;
        mem[1576] = 12'b001111001100;
        mem[1577] = 12'b001111001101;
        mem[1578] = 12'b001111001101;
        mem[1579] = 12'b001111001110;
        mem[1580] = 12'b001111001110;
        mem[1581] = 12'b001111001111;
        mem[1582] = 12'b001111010000;
        mem[1583] = 12'b001111010000;
        mem[1584] = 12'b001111010001;
        mem[1585] = 12'b001111010001;
        mem[1586] = 12'b001111010010;
        mem[1587] = 12'b001111010010;
        mem[1588] = 12'b001111010011;
        mem[1589] = 12'b001111010100;
        mem[1590] = 12'b001111010100;
        mem[1591] = 12'b001111010101;
        mem[1592] = 12'b001111010101;
        mem[1593] = 12'b001111010110;
        mem[1594] = 12'b001111010110;
        mem[1595] = 12'b001111010111;
        mem[1596] = 12'b001111010111;
        mem[1597] = 12'b001111011000;
        mem[1598] = 12'b001111011001;
        mem[1599] = 12'b001111011001;
        mem[1600] = 12'b001111011010;
        mem[1601] = 12'b001111011010;
        mem[1602] = 12'b001111011011;
        mem[1603] = 12'b001111011011;
        mem[1604] = 12'b001111011100;
        mem[1605] = 12'b001111011101;
        mem[1606] = 12'b001111011101;
        mem[1607] = 12'b001111011110;
        mem[1608] = 12'b001111011110;
        mem[1609] = 12'b001111011111;
        mem[1610] = 12'b001111011111;
        mem[1611] = 12'b001111100000;
        mem[1612] = 12'b001111100000;
        mem[1613] = 12'b001111100001;
        mem[1614] = 12'b001111100010;
        mem[1615] = 12'b001111100010;
        mem[1616] = 12'b001111100011;
        mem[1617] = 12'b001111100011;
        mem[1618] = 12'b001111100100;
        mem[1619] = 12'b001111100100;
        mem[1620] = 12'b001111100101;
        mem[1621] = 12'b001111100110;
        mem[1622] = 12'b001111100110;
        mem[1623] = 12'b001111100111;
        mem[1624] = 12'b001111100111;
        mem[1625] = 12'b001111101000;
        mem[1626] = 12'b001111101000;
        mem[1627] = 12'b001111101001;
        mem[1628] = 12'b001111101001;
        mem[1629] = 12'b001111101010;
        mem[1630] = 12'b001111101011;
        mem[1631] = 12'b001111101011;
        mem[1632] = 12'b001111101100;
        mem[1633] = 12'b001111101100;
        mem[1634] = 12'b001111101101;
        mem[1635] = 12'b001111101101;
        mem[1636] = 12'b001111101110;
        mem[1637] = 12'b001111101111;
        mem[1638] = 12'b001111101111;
        mem[1639] = 12'b001111110000;
        mem[1640] = 12'b001111110000;
        mem[1641] = 12'b001111110001;
        mem[1642] = 12'b001111110001;
        mem[1643] = 12'b001111110010;
        mem[1644] = 12'b001111110010;
        mem[1645] = 12'b001111110011;
        mem[1646] = 12'b001111110100;
        mem[1647] = 12'b001111110100;
        mem[1648] = 12'b001111110101;
        mem[1649] = 12'b001111110101;
        mem[1650] = 12'b001111110110;
        mem[1651] = 12'b001111110110;
        mem[1652] = 12'b001111110111;
        mem[1653] = 12'b001111110111;
        mem[1654] = 12'b001111111000;
        mem[1655] = 12'b001111111001;
        mem[1656] = 12'b001111111001;
        mem[1657] = 12'b001111111010;
        mem[1658] = 12'b001111111010;
        mem[1659] = 12'b001111111011;
        mem[1660] = 12'b001111111011;
        mem[1661] = 12'b001111111100;
        mem[1662] = 12'b001111111100;
        mem[1663] = 12'b001111111101;
        mem[1664] = 12'b001111111110;
        mem[1665] = 12'b001111111110;
        mem[1666] = 12'b001111111111;
        mem[1667] = 12'b001111111111;
        mem[1668] = 12'b010000000000;
        mem[1669] = 12'b010000000000;
        mem[1670] = 12'b010000000001;
        mem[1671] = 12'b010000000010;
        mem[1672] = 12'b010000000010;
        mem[1673] = 12'b010000000011;
        mem[1674] = 12'b010000000011;
        mem[1675] = 12'b010000000100;
        mem[1676] = 12'b010000000100;
        mem[1677] = 12'b010000000101;
        mem[1678] = 12'b010000000101;
        mem[1679] = 12'b010000000110;
        mem[1680] = 12'b010000000111;
        mem[1681] = 12'b010000000111;
        mem[1682] = 12'b010000001000;
        mem[1683] = 12'b010000001000;
        mem[1684] = 12'b010000001001;
        mem[1685] = 12'b010000001001;
        mem[1686] = 12'b010000001010;
        mem[1687] = 12'b010000001010;
        mem[1688] = 12'b010000001011;
        mem[1689] = 12'b010000001100;
        mem[1690] = 12'b010000001100;
        mem[1691] = 12'b010000001101;
        mem[1692] = 12'b010000001101;
        mem[1693] = 12'b010000001110;
        mem[1694] = 12'b010000001110;
        mem[1695] = 12'b010000001111;
        mem[1696] = 12'b010000001111;
        mem[1697] = 12'b010000010000;
        mem[1698] = 12'b010000010000;
        mem[1699] = 12'b010000010001;
        mem[1700] = 12'b010000010010;
        mem[1701] = 12'b010000010010;
        mem[1702] = 12'b010000010011;
        mem[1703] = 12'b010000010011;
        mem[1704] = 12'b010000010100;
        mem[1705] = 12'b010000010100;
        mem[1706] = 12'b010000010101;
        mem[1707] = 12'b010000010101;
        mem[1708] = 12'b010000010110;
        mem[1709] = 12'b010000010111;
        mem[1710] = 12'b010000010111;
        mem[1711] = 12'b010000011000;
        mem[1712] = 12'b010000011000;
        mem[1713] = 12'b010000011001;
        mem[1714] = 12'b010000011001;
        mem[1715] = 12'b010000011010;
        mem[1716] = 12'b010000011010;
        mem[1717] = 12'b010000011011;
        mem[1718] = 12'b010000011100;
        mem[1719] = 12'b010000011100;
        mem[1720] = 12'b010000011101;
        mem[1721] = 12'b010000011101;
        mem[1722] = 12'b010000011110;
        mem[1723] = 12'b010000011110;
        mem[1724] = 12'b010000011111;
        mem[1725] = 12'b010000011111;
        mem[1726] = 12'b010000100000;
        mem[1727] = 12'b010000100001;
        mem[1728] = 12'b010000100001;
        mem[1729] = 12'b010000100010;
        mem[1730] = 12'b010000100010;
        mem[1731] = 12'b010000100011;
        mem[1732] = 12'b010000100011;
        mem[1733] = 12'b010000100100;
        mem[1734] = 12'b010000100100;
        mem[1735] = 12'b010000100101;
        mem[1736] = 12'b010000100101;
        mem[1737] = 12'b010000100110;
        mem[1738] = 12'b010000100111;
        mem[1739] = 12'b010000100111;
        mem[1740] = 12'b010000101000;
        mem[1741] = 12'b010000101000;
        mem[1742] = 12'b010000101001;
        mem[1743] = 12'b010000101001;
        mem[1744] = 12'b010000101010;
        mem[1745] = 12'b010000101010;
        mem[1746] = 12'b010000101011;
        mem[1747] = 12'b010000101100;
        mem[1748] = 12'b010000101100;
        mem[1749] = 12'b010000101101;
        mem[1750] = 12'b010000101101;
        mem[1751] = 12'b010000101110;
        mem[1752] = 12'b010000101110;
        mem[1753] = 12'b010000101111;
        mem[1754] = 12'b010000101111;
        mem[1755] = 12'b010000110000;
        mem[1756] = 12'b010000110000;
        mem[1757] = 12'b010000110001;
        mem[1758] = 12'b010000110010;
        mem[1759] = 12'b010000110010;
        mem[1760] = 12'b010000110011;
        mem[1761] = 12'b010000110011;
        mem[1762] = 12'b010000110100;
        mem[1763] = 12'b010000110100;
        mem[1764] = 12'b010000110101;
        mem[1765] = 12'b010000110101;
        mem[1766] = 12'b010000110110;
        mem[1767] = 12'b010000110110;
        mem[1768] = 12'b010000110111;
        mem[1769] = 12'b010000111000;
        mem[1770] = 12'b010000111000;
        mem[1771] = 12'b010000111001;
        mem[1772] = 12'b010000111001;
        mem[1773] = 12'b010000111010;
        mem[1774] = 12'b010000111010;
        mem[1775] = 12'b010000111011;
        mem[1776] = 12'b010000111011;
        mem[1777] = 12'b010000111100;
        mem[1778] = 12'b010000111100;
        mem[1779] = 12'b010000111101;
        mem[1780] = 12'b010000111110;
        mem[1781] = 12'b010000111110;
        mem[1782] = 12'b010000111111;
        mem[1783] = 12'b010000111111;
        mem[1784] = 12'b010001000000;
        mem[1785] = 12'b010001000000;
        mem[1786] = 12'b010001000001;
        mem[1787] = 12'b010001000001;
        mem[1788] = 12'b010001000010;
        mem[1789] = 12'b010001000010;
        mem[1790] = 12'b010001000011;
        mem[1791] = 12'b010001000100;
        mem[1792] = 12'b010001000100;
        mem[1793] = 12'b010001000101;
        mem[1794] = 12'b010001000101;
        mem[1795] = 12'b010001000110;
        mem[1796] = 12'b010001000110;
        mem[1797] = 12'b010001000111;
        mem[1798] = 12'b010001000111;
        mem[1799] = 12'b010001001000;
        mem[1800] = 12'b010001001000;
        mem[1801] = 12'b010001001001;
        mem[1802] = 12'b010001001010;
        mem[1803] = 12'b010001001010;
        mem[1804] = 12'b010001001011;
        mem[1805] = 12'b010001001011;
        mem[1806] = 12'b010001001100;
        mem[1807] = 12'b010001001100;
        mem[1808] = 12'b010001001101;
        mem[1809] = 12'b010001001101;
        mem[1810] = 12'b010001001110;
        mem[1811] = 12'b010001001110;
        mem[1812] = 12'b010001001111;
        mem[1813] = 12'b010001001111;
        mem[1814] = 12'b010001010000;
        mem[1815] = 12'b010001010001;
        mem[1816] = 12'b010001010001;
        mem[1817] = 12'b010001010010;
        mem[1818] = 12'b010001010010;
        mem[1819] = 12'b010001010011;
        mem[1820] = 12'b010001010011;
        mem[1821] = 12'b010001010100;
        mem[1822] = 12'b010001010100;
        mem[1823] = 12'b010001010101;
        mem[1824] = 12'b010001010101;
        mem[1825] = 12'b010001010110;
        mem[1826] = 12'b010001010111;
        mem[1827] = 12'b010001010111;
        mem[1828] = 12'b010001011000;
        mem[1829] = 12'b010001011000;
        mem[1830] = 12'b010001011001;
        mem[1831] = 12'b010001011001;
        mem[1832] = 12'b010001011010;
        mem[1833] = 12'b010001011010;
        mem[1834] = 12'b010001011011;
        mem[1835] = 12'b010001011011;
        mem[1836] = 12'b010001011100;
        mem[1837] = 12'b010001011100;
        mem[1838] = 12'b010001011101;
        mem[1839] = 12'b010001011110;
        mem[1840] = 12'b010001011110;
        mem[1841] = 12'b010001011111;
        mem[1842] = 12'b010001011111;
        mem[1843] = 12'b010001100000;
        mem[1844] = 12'b010001100000;
        mem[1845] = 12'b010001100001;
        mem[1846] = 12'b010001100001;
        mem[1847] = 12'b010001100010;
        mem[1848] = 12'b010001100010;
        mem[1849] = 12'b010001100011;
        mem[1850] = 12'b010001100011;
        mem[1851] = 12'b010001100100;
        mem[1852] = 12'b010001100101;
        mem[1853] = 12'b010001100101;
        mem[1854] = 12'b010001100110;
        mem[1855] = 12'b010001100110;
        mem[1856] = 12'b010001100111;
        mem[1857] = 12'b010001100111;
        mem[1858] = 12'b010001101000;
        mem[1859] = 12'b010001101000;
        mem[1860] = 12'b010001101001;
        mem[1861] = 12'b010001101001;
        mem[1862] = 12'b010001101010;
        mem[1863] = 12'b010001101010;
        mem[1864] = 12'b010001101011;
        mem[1865] = 12'b010001101011;
        mem[1866] = 12'b010001101100;
        mem[1867] = 12'b010001101101;
        mem[1868] = 12'b010001101101;
        mem[1869] = 12'b010001101110;
        mem[1870] = 12'b010001101110;
        mem[1871] = 12'b010001101111;
        mem[1872] = 12'b010001101111;
        mem[1873] = 12'b010001110000;
        mem[1874] = 12'b010001110000;
        mem[1875] = 12'b010001110001;
        mem[1876] = 12'b010001110001;
        mem[1877] = 12'b010001110010;
        mem[1878] = 12'b010001110010;
        mem[1879] = 12'b010001110011;
        mem[1880] = 12'b010001110100;
        mem[1881] = 12'b010001110100;
        mem[1882] = 12'b010001110101;
        mem[1883] = 12'b010001110101;
        mem[1884] = 12'b010001110110;
        mem[1885] = 12'b010001110110;
        mem[1886] = 12'b010001110111;
        mem[1887] = 12'b010001110111;
        mem[1888] = 12'b010001111000;
        mem[1889] = 12'b010001111000;
        mem[1890] = 12'b010001111001;
        mem[1891] = 12'b010001111001;
        mem[1892] = 12'b010001111010;
        mem[1893] = 12'b010001111010;
        mem[1894] = 12'b010001111011;
        mem[1895] = 12'b010001111100;
        mem[1896] = 12'b010001111100;
        mem[1897] = 12'b010001111101;
        mem[1898] = 12'b010001111101;
        mem[1899] = 12'b010001111110;
        mem[1900] = 12'b010001111110;
        mem[1901] = 12'b010001111111;
        mem[1902] = 12'b010001111111;
        mem[1903] = 12'b010010000000;
        mem[1904] = 12'b010010000000;
        mem[1905] = 12'b010010000001;
        mem[1906] = 12'b010010000001;
        mem[1907] = 12'b010010000010;
        mem[1908] = 12'b010010000010;
        mem[1909] = 12'b010010000011;
        mem[1910] = 12'b010010000011;
        mem[1911] = 12'b010010000100;
        mem[1912] = 12'b010010000101;
        mem[1913] = 12'b010010000101;
        mem[1914] = 12'b010010000110;
        mem[1915] = 12'b010010000110;
        mem[1916] = 12'b010010000111;
        mem[1917] = 12'b010010000111;
        mem[1918] = 12'b010010001000;
        mem[1919] = 12'b010010001000;
        mem[1920] = 12'b010010001001;
        mem[1921] = 12'b010010001001;
        mem[1922] = 12'b010010001010;
        mem[1923] = 12'b010010001010;
        mem[1924] = 12'b010010001011;
        mem[1925] = 12'b010010001011;
        mem[1926] = 12'b010010001100;
        mem[1927] = 12'b010010001101;
        mem[1928] = 12'b010010001101;
        mem[1929] = 12'b010010001110;
        mem[1930] = 12'b010010001110;
        mem[1931] = 12'b010010001111;
        mem[1932] = 12'b010010001111;
        mem[1933] = 12'b010010010000;
        mem[1934] = 12'b010010010000;
        mem[1935] = 12'b010010010001;
        mem[1936] = 12'b010010010001;
        mem[1937] = 12'b010010010010;
        mem[1938] = 12'b010010010010;
        mem[1939] = 12'b010010010011;
        mem[1940] = 12'b010010010011;
        mem[1941] = 12'b010010010100;
        mem[1942] = 12'b010010010100;
        mem[1943] = 12'b010010010101;
        mem[1944] = 12'b010010010101;
        mem[1945] = 12'b010010010110;
        mem[1946] = 12'b010010010111;
        mem[1947] = 12'b010010010111;
        mem[1948] = 12'b010010011000;
        mem[1949] = 12'b010010011000;
        mem[1950] = 12'b010010011001;
        mem[1951] = 12'b010010011001;
        mem[1952] = 12'b010010011010;
        mem[1953] = 12'b010010011010;
        mem[1954] = 12'b010010011011;
        mem[1955] = 12'b010010011011;
        mem[1956] = 12'b010010011100;
        mem[1957] = 12'b010010011100;
        mem[1958] = 12'b010010011101;
        mem[1959] = 12'b010010011101;
        mem[1960] = 12'b010010011110;
        mem[1961] = 12'b010010011110;
        mem[1962] = 12'b010010011111;
        mem[1963] = 12'b010010011111;
        mem[1964] = 12'b010010100000;
        mem[1965] = 12'b010010100001;
        mem[1966] = 12'b010010100001;
        mem[1967] = 12'b010010100010;
        mem[1968] = 12'b010010100010;
        mem[1969] = 12'b010010100011;
        mem[1970] = 12'b010010100011;
        mem[1971] = 12'b010010100100;
        mem[1972] = 12'b010010100100;
        mem[1973] = 12'b010010100101;
        mem[1974] = 12'b010010100101;
        mem[1975] = 12'b010010100110;
        mem[1976] = 12'b010010100110;
        mem[1977] = 12'b010010100111;
        mem[1978] = 12'b010010100111;
        mem[1979] = 12'b010010101000;
        mem[1980] = 12'b010010101000;
        mem[1981] = 12'b010010101001;
        mem[1982] = 12'b010010101001;
        mem[1983] = 12'b010010101010;
        mem[1984] = 12'b010010101010;
        mem[1985] = 12'b010010101011;
        mem[1986] = 12'b010010101100;
        mem[1987] = 12'b010010101100;
        mem[1988] = 12'b010010101101;
        mem[1989] = 12'b010010101101;
        mem[1990] = 12'b010010101110;
        mem[1991] = 12'b010010101110;
        mem[1992] = 12'b010010101111;
        mem[1993] = 12'b010010101111;
        mem[1994] = 12'b010010110000;
        mem[1995] = 12'b010010110000;
        mem[1996] = 12'b010010110001;
        mem[1997] = 12'b010010110001;
        mem[1998] = 12'b010010110010;
        mem[1999] = 12'b010010110010;
        mem[2000] = 12'b010010110011;
        mem[2001] = 12'b010010110011;
        mem[2002] = 12'b010010110100;
        mem[2003] = 12'b010010110100;
        mem[2004] = 12'b010010110101;
        mem[2005] = 12'b010010110101;
        mem[2006] = 12'b010010110110;
        mem[2007] = 12'b010010110110;
        mem[2008] = 12'b010010110111;
        mem[2009] = 12'b010010110111;
        mem[2010] = 12'b010010111000;
        mem[2011] = 12'b010010111001;
        mem[2012] = 12'b010010111001;
        mem[2013] = 12'b010010111010;
        mem[2014] = 12'b010010111010;
        mem[2015] = 12'b010010111011;
        mem[2016] = 12'b010010111011;
        mem[2017] = 12'b010010111100;
        mem[2018] = 12'b010010111100;
        mem[2019] = 12'b010010111101;
        mem[2020] = 12'b010010111101;
        mem[2021] = 12'b010010111110;
        mem[2022] = 12'b010010111110;
        mem[2023] = 12'b010010111111;
        mem[2024] = 12'b010010111111;
        mem[2025] = 12'b010011000000;
        mem[2026] = 12'b010011000000;
        mem[2027] = 12'b010011000001;
        mem[2028] = 12'b010011000001;
        mem[2029] = 12'b010011000010;
        mem[2030] = 12'b010011000010;
        mem[2031] = 12'b010011000011;
        mem[2032] = 12'b010011000011;
        mem[2033] = 12'b010011000100;
        mem[2034] = 12'b010011000100;
        mem[2035] = 12'b010011000101;
        mem[2036] = 12'b010011000101;
        mem[2037] = 12'b010011000110;
        mem[2038] = 12'b010011000110;
        mem[2039] = 12'b010011000111;
        mem[2040] = 12'b010011001000;
        mem[2041] = 12'b010011001000;
        mem[2042] = 12'b010011001001;
        mem[2043] = 12'b010011001001;
        mem[2044] = 12'b010011001010;
        mem[2045] = 12'b010011001010;
        mem[2046] = 12'b010011001011;
        mem[2047] = 12'b010011001011;
        mem[2048] = 12'b010011001100;
        mem[2049] = 12'b010011001100;
        mem[2050] = 12'b010011001101;
        mem[2051] = 12'b010011001101;
        mem[2052] = 12'b010011001110;
        mem[2053] = 12'b010011001110;
        mem[2054] = 12'b010011001111;
        mem[2055] = 12'b010011001111;
        mem[2056] = 12'b010011010000;
        mem[2057] = 12'b010011010000;
        mem[2058] = 12'b010011010001;
        mem[2059] = 12'b010011010001;
        mem[2060] = 12'b010011010010;
        mem[2061] = 12'b010011010010;
        mem[2062] = 12'b010011010011;
        mem[2063] = 12'b010011010011;
        mem[2064] = 12'b010011010100;
        mem[2065] = 12'b010011010100;
        mem[2066] = 12'b010011010101;
        mem[2067] = 12'b010011010101;
        mem[2068] = 12'b010011010110;
        mem[2069] = 12'b010011010110;
        mem[2070] = 12'b010011010111;
        mem[2071] = 12'b010011010111;
        mem[2072] = 12'b010011011000;
        mem[2073] = 12'b010011011000;
        mem[2074] = 12'b010011011001;
        mem[2075] = 12'b010011011001;
        mem[2076] = 12'b010011011010;
        mem[2077] = 12'b010011011011;
        mem[2078] = 12'b010011011011;
        mem[2079] = 12'b010011011100;
        mem[2080] = 12'b010011011100;
        mem[2081] = 12'b010011011101;
        mem[2082] = 12'b010011011101;
        mem[2083] = 12'b010011011110;
        mem[2084] = 12'b010011011110;
        mem[2085] = 12'b010011011111;
        mem[2086] = 12'b010011011111;
        mem[2087] = 12'b010011100000;
        mem[2088] = 12'b010011100000;
        mem[2089] = 12'b010011100001;
        mem[2090] = 12'b010011100001;
        mem[2091] = 12'b010011100010;
        mem[2092] = 12'b010011100010;
        mem[2093] = 12'b010011100011;
        mem[2094] = 12'b010011100011;
        mem[2095] = 12'b010011100100;
        mem[2096] = 12'b010011100100;
        mem[2097] = 12'b010011100101;
        mem[2098] = 12'b010011100101;
        mem[2099] = 12'b010011100110;
        mem[2100] = 12'b010011100110;
        mem[2101] = 12'b010011100111;
        mem[2102] = 12'b010011100111;
        mem[2103] = 12'b010011101000;
        mem[2104] = 12'b010011101000;
        mem[2105] = 12'b010011101001;
        mem[2106] = 12'b010011101001;
        mem[2107] = 12'b010011101010;
        mem[2108] = 12'b010011101010;
        mem[2109] = 12'b010011101011;
        mem[2110] = 12'b010011101011;
        mem[2111] = 12'b010011101100;
        mem[2112] = 12'b010011101100;
        mem[2113] = 12'b010011101101;
        mem[2114] = 12'b010011101101;
        mem[2115] = 12'b010011101110;
        mem[2116] = 12'b010011101110;
        mem[2117] = 12'b010011101111;
        mem[2118] = 12'b010011101111;
        mem[2119] = 12'b010011110000;
        mem[2120] = 12'b010011110000;
        mem[2121] = 12'b010011110001;
        mem[2122] = 12'b010011110001;
        mem[2123] = 12'b010011110010;
        mem[2124] = 12'b010011110010;
        mem[2125] = 12'b010011110011;
        mem[2126] = 12'b010011110011;
        mem[2127] = 12'b010011110100;
        mem[2128] = 12'b010011110100;
        mem[2129] = 12'b010011110101;
        mem[2130] = 12'b010011110101;
        mem[2131] = 12'b010011110110;
        mem[2132] = 12'b010011110110;
        mem[2133] = 12'b010011110111;
        mem[2134] = 12'b010011110111;
        mem[2135] = 12'b010011111000;
        mem[2136] = 12'b010011111000;
        mem[2137] = 12'b010011111001;
        mem[2138] = 12'b010011111001;
        mem[2139] = 12'b010011111010;
        mem[2140] = 12'b010011111010;
        mem[2141] = 12'b010011111011;
        mem[2142] = 12'b010011111011;
        mem[2143] = 12'b010011111100;
        mem[2144] = 12'b010011111100;
        mem[2145] = 12'b010011111101;
        mem[2146] = 12'b010011111101;
        mem[2147] = 12'b010011111110;
        mem[2148] = 12'b010011111110;
        mem[2149] = 12'b010011111111;
        mem[2150] = 12'b010011111111;
        mem[2151] = 12'b010100000000;
        mem[2152] = 12'b010100000000;
        mem[2153] = 12'b010100000001;
        mem[2154] = 12'b010100000001;
        mem[2155] = 12'b010100000010;
        mem[2156] = 12'b010100000010;
        mem[2157] = 12'b010100000011;
        mem[2158] = 12'b010100000011;
        mem[2159] = 12'b010100000100;
        mem[2160] = 12'b010100000100;
        mem[2161] = 12'b010100000101;
        mem[2162] = 12'b010100000101;
        mem[2163] = 12'b010100000110;
        mem[2164] = 12'b010100000110;
        mem[2165] = 12'b010100000111;
        mem[2166] = 12'b010100000111;
        mem[2167] = 12'b010100001000;
        mem[2168] = 12'b010100001000;
        mem[2169] = 12'b010100001001;
        mem[2170] = 12'b010100001001;
        mem[2171] = 12'b010100001010;
        mem[2172] = 12'b010100001010;
        mem[2173] = 12'b010100001011;
        mem[2174] = 12'b010100001011;
        mem[2175] = 12'b010100001100;
        mem[2176] = 12'b010100001100;
        mem[2177] = 12'b010100001101;
        mem[2178] = 12'b010100001101;
        mem[2179] = 12'b010100001110;
        mem[2180] = 12'b010100001110;
        mem[2181] = 12'b010100001111;
        mem[2182] = 12'b010100001111;
        mem[2183] = 12'b010100010000;
        mem[2184] = 12'b010100010000;
        mem[2185] = 12'b010100010001;
        mem[2186] = 12'b010100010001;
        mem[2187] = 12'b010100010010;
        mem[2188] = 12'b010100010010;
        mem[2189] = 12'b010100010011;
        mem[2190] = 12'b010100010011;
        mem[2191] = 12'b010100010100;
        mem[2192] = 12'b010100010100;
        mem[2193] = 12'b010100010101;
        mem[2194] = 12'b010100010101;
        mem[2195] = 12'b010100010110;
        mem[2196] = 12'b010100010110;
        mem[2197] = 12'b010100010111;
        mem[2198] = 12'b010100010111;
        mem[2199] = 12'b010100011000;
        mem[2200] = 12'b010100011000;
        mem[2201] = 12'b010100011001;
        mem[2202] = 12'b010100011001;
        mem[2203] = 12'b010100011010;
        mem[2204] = 12'b010100011010;
        mem[2205] = 12'b010100011011;
        mem[2206] = 12'b010100011011;
        mem[2207] = 12'b010100011100;
        mem[2208] = 12'b010100011100;
        mem[2209] = 12'b010100011101;
        mem[2210] = 12'b010100011101;
        mem[2211] = 12'b010100011110;
        mem[2212] = 12'b010100011110;
        mem[2213] = 12'b010100011111;
        mem[2214] = 12'b010100011111;
        mem[2215] = 12'b010100100000;
        mem[2216] = 12'b010100100000;
        mem[2217] = 12'b010100100001;
        mem[2218] = 12'b010100100001;
        mem[2219] = 12'b010100100010;
        mem[2220] = 12'b010100100010;
        mem[2221] = 12'b010100100011;
        mem[2222] = 12'b010100100011;
        mem[2223] = 12'b010100100100;
        mem[2224] = 12'b010100100100;
        mem[2225] = 12'b010100100101;
        mem[2226] = 12'b010100100101;
        mem[2227] = 12'b010100100110;
        mem[2228] = 12'b010100100110;
        mem[2229] = 12'b010100100111;
        mem[2230] = 12'b010100100111;
        mem[2231] = 12'b010100101000;
        mem[2232] = 12'b010100101000;
        mem[2233] = 12'b010100101001;
        mem[2234] = 12'b010100101001;
        mem[2235] = 12'b010100101010;
        mem[2236] = 12'b010100101010;
        mem[2237] = 12'b010100101011;
        mem[2238] = 12'b010100101011;
        mem[2239] = 12'b010100101100;
        mem[2240] = 12'b010100101100;
        mem[2241] = 12'b010100101101;
        mem[2242] = 12'b010100101101;
        mem[2243] = 12'b010100101110;
        mem[2244] = 12'b010100101110;
        mem[2245] = 12'b010100101111;
        mem[2246] = 12'b010100101111;
        mem[2247] = 12'b010100110000;
        mem[2248] = 12'b010100110000;
        mem[2249] = 12'b010100110001;
        mem[2250] = 12'b010100110001;
        mem[2251] = 12'b010100110010;
        mem[2252] = 12'b010100110010;
        mem[2253] = 12'b010100110010;
        mem[2254] = 12'b010100110011;
        mem[2255] = 12'b010100110011;
        mem[2256] = 12'b010100110100;
        mem[2257] = 12'b010100110100;
        mem[2258] = 12'b010100110101;
        mem[2259] = 12'b010100110101;
        mem[2260] = 12'b010100110110;
        mem[2261] = 12'b010100110110;
        mem[2262] = 12'b010100110111;
        mem[2263] = 12'b010100110111;
        mem[2264] = 12'b010100111000;
        mem[2265] = 12'b010100111000;
        mem[2266] = 12'b010100111001;
        mem[2267] = 12'b010100111001;
        mem[2268] = 12'b010100111010;
        mem[2269] = 12'b010100111010;
        mem[2270] = 12'b010100111011;
        mem[2271] = 12'b010100111011;
        mem[2272] = 12'b010100111100;
        mem[2273] = 12'b010100111100;
        mem[2274] = 12'b010100111101;
        mem[2275] = 12'b010100111101;
        mem[2276] = 12'b010100111110;
        mem[2277] = 12'b010100111110;
        mem[2278] = 12'b010100111111;
        mem[2279] = 12'b010100111111;
        mem[2280] = 12'b010101000000;
        mem[2281] = 12'b010101000000;
        mem[2282] = 12'b010101000001;
        mem[2283] = 12'b010101000001;
        mem[2284] = 12'b010101000010;
        mem[2285] = 12'b010101000010;
        mem[2286] = 12'b010101000011;
        mem[2287] = 12'b010101000011;
        mem[2288] = 12'b010101000100;
        mem[2289] = 12'b010101000100;
        mem[2290] = 12'b010101000100;
        mem[2291] = 12'b010101000101;
        mem[2292] = 12'b010101000101;
        mem[2293] = 12'b010101000110;
        mem[2294] = 12'b010101000110;
        mem[2295] = 12'b010101000111;
        mem[2296] = 12'b010101000111;
        mem[2297] = 12'b010101001000;
        mem[2298] = 12'b010101001000;
        mem[2299] = 12'b010101001001;
        mem[2300] = 12'b010101001001;
        mem[2301] = 12'b010101001010;
        mem[2302] = 12'b010101001010;
        mem[2303] = 12'b010101001011;
        mem[2304] = 12'b010101001011;
        mem[2305] = 12'b010101001100;
        mem[2306] = 12'b010101001100;
        mem[2307] = 12'b010101001101;
        mem[2308] = 12'b010101001101;
        mem[2309] = 12'b010101001110;
        mem[2310] = 12'b010101001110;
        mem[2311] = 12'b010101001111;
        mem[2312] = 12'b010101001111;
        mem[2313] = 12'b010101010000;
        mem[2314] = 12'b010101010000;
        mem[2315] = 12'b010101010001;
        mem[2316] = 12'b010101010001;
        mem[2317] = 12'b010101010001;
        mem[2318] = 12'b010101010010;
        mem[2319] = 12'b010101010010;
        mem[2320] = 12'b010101010011;
        mem[2321] = 12'b010101010011;
        mem[2322] = 12'b010101010100;
        mem[2323] = 12'b010101010100;
        mem[2324] = 12'b010101010101;
        mem[2325] = 12'b010101010101;
        mem[2326] = 12'b010101010110;
        mem[2327] = 12'b010101010110;
        mem[2328] = 12'b010101010111;
        mem[2329] = 12'b010101010111;
        mem[2330] = 12'b010101011000;
        mem[2331] = 12'b010101011000;
        mem[2332] = 12'b010101011001;
        mem[2333] = 12'b010101011001;
        mem[2334] = 12'b010101011010;
        mem[2335] = 12'b010101011010;
        mem[2336] = 12'b010101011011;
        mem[2337] = 12'b010101011011;
        mem[2338] = 12'b010101011100;
        mem[2339] = 12'b010101011100;
        mem[2340] = 12'b010101011101;
        mem[2341] = 12'b010101011101;
        mem[2342] = 12'b010101011101;
        mem[2343] = 12'b010101011110;
        mem[2344] = 12'b010101011110;
        mem[2345] = 12'b010101011111;
        mem[2346] = 12'b010101011111;
        mem[2347] = 12'b010101100000;
        mem[2348] = 12'b010101100000;
        mem[2349] = 12'b010101100001;
        mem[2350] = 12'b010101100001;
        mem[2351] = 12'b010101100010;
        mem[2352] = 12'b010101100010;
        mem[2353] = 12'b010101100011;
        mem[2354] = 12'b010101100011;
        mem[2355] = 12'b010101100100;
        mem[2356] = 12'b010101100100;
        mem[2357] = 12'b010101100101;
        mem[2358] = 12'b010101100101;
        mem[2359] = 12'b010101100110;
        mem[2360] = 12'b010101100110;
        mem[2361] = 12'b010101100110;
        mem[2362] = 12'b010101100111;
        mem[2363] = 12'b010101100111;
        mem[2364] = 12'b010101101000;
        mem[2365] = 12'b010101101000;
        mem[2366] = 12'b010101101001;
        mem[2367] = 12'b010101101001;
        mem[2368] = 12'b010101101010;
        mem[2369] = 12'b010101101010;
        mem[2370] = 12'b010101101011;
        mem[2371] = 12'b010101101011;
        mem[2372] = 12'b010101101100;
        mem[2373] = 12'b010101101100;
        mem[2374] = 12'b010101101101;
        mem[2375] = 12'b010101101101;
        mem[2376] = 12'b010101101110;
        mem[2377] = 12'b010101101110;
        mem[2378] = 12'b010101101111;
        mem[2379] = 12'b010101101111;
        mem[2380] = 12'b010101101111;
        mem[2381] = 12'b010101110000;
        mem[2382] = 12'b010101110000;
        mem[2383] = 12'b010101110001;
        mem[2384] = 12'b010101110001;
        mem[2385] = 12'b010101110010;
        mem[2386] = 12'b010101110010;
        mem[2387] = 12'b010101110011;
        mem[2388] = 12'b010101110011;
        mem[2389] = 12'b010101110100;
        mem[2390] = 12'b010101110100;
        mem[2391] = 12'b010101110101;
        mem[2392] = 12'b010101110101;
        mem[2393] = 12'b010101110110;
        mem[2394] = 12'b010101110110;
        mem[2395] = 12'b010101110111;
        mem[2396] = 12'b010101110111;
        mem[2397] = 12'b010101110111;
        mem[2398] = 12'b010101111000;
        mem[2399] = 12'b010101111000;
        mem[2400] = 12'b010101111001;
        mem[2401] = 12'b010101111001;
        mem[2402] = 12'b010101111010;
        mem[2403] = 12'b010101111010;
        mem[2404] = 12'b010101111011;
        mem[2405] = 12'b010101111011;
        mem[2406] = 12'b010101111100;
        mem[2407] = 12'b010101111100;
        mem[2408] = 12'b010101111101;
        mem[2409] = 12'b010101111101;
        mem[2410] = 12'b010101111110;
        mem[2411] = 12'b010101111110;
        mem[2412] = 12'b010101111110;
        mem[2413] = 12'b010101111111;
        mem[2414] = 12'b010101111111;
        mem[2415] = 12'b010110000000;
        mem[2416] = 12'b010110000000;
        mem[2417] = 12'b010110000001;
        mem[2418] = 12'b010110000001;
        mem[2419] = 12'b010110000010;
        mem[2420] = 12'b010110000010;
        mem[2421] = 12'b010110000011;
        mem[2422] = 12'b010110000011;
        mem[2423] = 12'b010110000100;
        mem[2424] = 12'b010110000100;
        mem[2425] = 12'b010110000101;
        mem[2426] = 12'b010110000101;
        mem[2427] = 12'b010110000101;
        mem[2428] = 12'b010110000110;
        mem[2429] = 12'b010110000110;
        mem[2430] = 12'b010110000111;
        mem[2431] = 12'b010110000111;
        mem[2432] = 12'b010110001000;
        mem[2433] = 12'b010110001000;
        mem[2434] = 12'b010110001001;
        mem[2435] = 12'b010110001001;
        mem[2436] = 12'b010110001010;
        mem[2437] = 12'b010110001010;
        mem[2438] = 12'b010110001011;
        mem[2439] = 12'b010110001011;
        mem[2440] = 12'b010110001100;
        mem[2441] = 12'b010110001100;
        mem[2442] = 12'b010110001100;
        mem[2443] = 12'b010110001101;
        mem[2444] = 12'b010110001101;
        mem[2445] = 12'b010110001110;
        mem[2446] = 12'b010110001110;
        mem[2447] = 12'b010110001111;
        mem[2448] = 12'b010110001111;
        mem[2449] = 12'b010110010000;
        mem[2450] = 12'b010110010000;
        mem[2451] = 12'b010110010001;
        mem[2452] = 12'b010110010001;
        mem[2453] = 12'b010110010010;
        mem[2454] = 12'b010110010010;
        mem[2455] = 12'b010110010010;
        mem[2456] = 12'b010110010011;
        mem[2457] = 12'b010110010011;
        mem[2458] = 12'b010110010100;
        mem[2459] = 12'b010110010100;
        mem[2460] = 12'b010110010101;
        mem[2461] = 12'b010110010101;
        mem[2462] = 12'b010110010110;
        mem[2463] = 12'b010110010110;
        mem[2464] = 12'b010110010111;
        mem[2465] = 12'b010110010111;
        mem[2466] = 12'b010110011000;
        mem[2467] = 12'b010110011000;
        mem[2468] = 12'b010110011000;
        mem[2469] = 12'b010110011001;
        mem[2470] = 12'b010110011001;
        mem[2471] = 12'b010110011010;
        mem[2472] = 12'b010110011010;
        mem[2473] = 12'b010110011011;
        mem[2474] = 12'b010110011011;
        mem[2475] = 12'b010110011100;
        mem[2476] = 12'b010110011100;
        mem[2477] = 12'b010110011101;
        mem[2478] = 12'b010110011101;
        mem[2479] = 12'b010110011101;
        mem[2480] = 12'b010110011110;
        mem[2481] = 12'b010110011110;
        mem[2482] = 12'b010110011111;
        mem[2483] = 12'b010110011111;
        mem[2484] = 12'b010110100000;
        mem[2485] = 12'b010110100000;
        mem[2486] = 12'b010110100001;
        mem[2487] = 12'b010110100001;
        mem[2488] = 12'b010110100010;
        mem[2489] = 12'b010110100010;
        mem[2490] = 12'b010110100011;
        mem[2491] = 12'b010110100011;
        mem[2492] = 12'b010110100011;
        mem[2493] = 12'b010110100100;
        mem[2494] = 12'b010110100100;
        mem[2495] = 12'b010110100101;
        mem[2496] = 12'b010110100101;
        mem[2497] = 12'b010110100110;
        mem[2498] = 12'b010110100110;
        mem[2499] = 12'b010110100111;
        mem[2500] = 12'b010110100111;
        mem[2501] = 12'b010110101000;
        mem[2502] = 12'b010110101000;
        mem[2503] = 12'b010110101000;
        mem[2504] = 12'b010110101001;
        mem[2505] = 12'b010110101001;
        mem[2506] = 12'b010110101010;
        mem[2507] = 12'b010110101010;
        mem[2508] = 12'b010110101011;
        mem[2509] = 12'b010110101011;
        mem[2510] = 12'b010110101100;
        mem[2511] = 12'b010110101100;
        mem[2512] = 12'b010110101101;
        mem[2513] = 12'b010110101101;
        mem[2514] = 12'b010110101101;
        mem[2515] = 12'b010110101110;
        mem[2516] = 12'b010110101110;
        mem[2517] = 12'b010110101111;
        mem[2518] = 12'b010110101111;
        mem[2519] = 12'b010110110000;
        mem[2520] = 12'b010110110000;
        mem[2521] = 12'b010110110001;
        mem[2522] = 12'b010110110001;
        mem[2523] = 12'b010110110001;
        mem[2524] = 12'b010110110010;
        mem[2525] = 12'b010110110010;
        mem[2526] = 12'b010110110011;
        mem[2527] = 12'b010110110011;
        mem[2528] = 12'b010110110100;
        mem[2529] = 12'b010110110100;
        mem[2530] = 12'b010110110101;
        mem[2531] = 12'b010110110101;
        mem[2532] = 12'b010110110110;
        mem[2533] = 12'b010110110110;
        mem[2534] = 12'b010110110110;
        mem[2535] = 12'b010110110111;
        mem[2536] = 12'b010110110111;
        mem[2537] = 12'b010110111000;
        mem[2538] = 12'b010110111000;
        mem[2539] = 12'b010110111001;
        mem[2540] = 12'b010110111001;
        mem[2541] = 12'b010110111010;
        mem[2542] = 12'b010110111010;
        mem[2543] = 12'b010110111010;
        mem[2544] = 12'b010110111011;
        mem[2545] = 12'b010110111011;
        mem[2546] = 12'b010110111100;
        mem[2547] = 12'b010110111100;
        mem[2548] = 12'b010110111101;
        mem[2549] = 12'b010110111101;
        mem[2550] = 12'b010110111110;
        mem[2551] = 12'b010110111110;
        mem[2552] = 12'b010110111111;
        mem[2553] = 12'b010110111111;
        mem[2554] = 12'b010110111111;
        mem[2555] = 12'b010111000000;
        mem[2556] = 12'b010111000000;
        mem[2557] = 12'b010111000001;
        mem[2558] = 12'b010111000001;
        mem[2559] = 12'b010111000010;
        mem[2560] = 12'b010111000010;
        mem[2561] = 12'b010111000011;
        mem[2562] = 12'b010111000011;
        mem[2563] = 12'b010111000011;
        mem[2564] = 12'b010111000100;
        mem[2565] = 12'b010111000100;
        mem[2566] = 12'b010111000101;
        mem[2567] = 12'b010111000101;
        mem[2568] = 12'b010111000110;
        mem[2569] = 12'b010111000110;
        mem[2570] = 12'b010111000111;
        mem[2571] = 12'b010111000111;
        mem[2572] = 12'b010111000111;
        mem[2573] = 12'b010111001000;
        mem[2574] = 12'b010111001000;
        mem[2575] = 12'b010111001001;
        mem[2576] = 12'b010111001001;
        mem[2577] = 12'b010111001010;
        mem[2578] = 12'b010111001010;
        mem[2579] = 12'b010111001011;
        mem[2580] = 12'b010111001011;
        mem[2581] = 12'b010111001011;
        mem[2582] = 12'b010111001100;
        mem[2583] = 12'b010111001100;
        mem[2584] = 12'b010111001101;
        mem[2585] = 12'b010111001101;
        mem[2586] = 12'b010111001110;
        mem[2587] = 12'b010111001110;
        mem[2588] = 12'b010111001111;
        mem[2589] = 12'b010111001111;
        mem[2590] = 12'b010111001111;
        mem[2591] = 12'b010111010000;
        mem[2592] = 12'b010111010000;
        mem[2593] = 12'b010111010001;
        mem[2594] = 12'b010111010001;
        mem[2595] = 12'b010111010010;
        mem[2596] = 12'b010111010010;
        mem[2597] = 12'b010111010010;
        mem[2598] = 12'b010111010011;
        mem[2599] = 12'b010111010011;
        mem[2600] = 12'b010111010100;
        mem[2601] = 12'b010111010100;
        mem[2602] = 12'b010111010101;
        mem[2603] = 12'b010111010101;
        mem[2604] = 12'b010111010110;
        mem[2605] = 12'b010111010110;
        mem[2606] = 12'b010111010110;
        mem[2607] = 12'b010111010111;
        mem[2608] = 12'b010111010111;
        mem[2609] = 12'b010111011000;
        mem[2610] = 12'b010111011000;
        mem[2611] = 12'b010111011001;
        mem[2612] = 12'b010111011001;
        mem[2613] = 12'b010111011010;
        mem[2614] = 12'b010111011010;
        mem[2615] = 12'b010111011010;
        mem[2616] = 12'b010111011011;
        mem[2617] = 12'b010111011011;
        mem[2618] = 12'b010111011100;
        mem[2619] = 12'b010111011100;
        mem[2620] = 12'b010111011101;
        mem[2621] = 12'b010111011101;
        mem[2622] = 12'b010111011101;
        mem[2623] = 12'b010111011110;
        mem[2624] = 12'b010111011110;
        mem[2625] = 12'b010111011111;
        mem[2626] = 12'b010111011111;
        mem[2627] = 12'b010111100000;
        mem[2628] = 12'b010111100000;
        mem[2629] = 12'b010111100001;
        mem[2630] = 12'b010111100001;
        mem[2631] = 12'b010111100001;
        mem[2632] = 12'b010111100010;
        mem[2633] = 12'b010111100010;
        mem[2634] = 12'b010111100011;
        mem[2635] = 12'b010111100011;
        mem[2636] = 12'b010111100100;
        mem[2637] = 12'b010111100100;
        mem[2638] = 12'b010111100100;
        mem[2639] = 12'b010111100101;
        mem[2640] = 12'b010111100101;
        mem[2641] = 12'b010111100110;
        mem[2642] = 12'b010111100110;
        mem[2643] = 12'b010111100111;
        mem[2644] = 12'b010111100111;
        mem[2645] = 12'b010111100111;
        mem[2646] = 12'b010111101000;
        mem[2647] = 12'b010111101000;
        mem[2648] = 12'b010111101001;
        mem[2649] = 12'b010111101001;
        mem[2650] = 12'b010111101010;
        mem[2651] = 12'b010111101010;
        mem[2652] = 12'b010111101011;
        mem[2653] = 12'b010111101011;
        mem[2654] = 12'b010111101011;
        mem[2655] = 12'b010111101100;
        mem[2656] = 12'b010111101100;
        mem[2657] = 12'b010111101101;
        mem[2658] = 12'b010111101101;
        mem[2659] = 12'b010111101110;
        mem[2660] = 12'b010111101110;
        mem[2661] = 12'b010111101110;
        mem[2662] = 12'b010111101111;
        mem[2663] = 12'b010111101111;
        mem[2664] = 12'b010111110000;
        mem[2665] = 12'b010111110000;
        mem[2666] = 12'b010111110001;
        mem[2667] = 12'b010111110001;
        mem[2668] = 12'b010111110001;
        mem[2669] = 12'b010111110010;
        mem[2670] = 12'b010111110010;
        mem[2671] = 12'b010111110011;
        mem[2672] = 12'b010111110011;
        mem[2673] = 12'b010111110100;
        mem[2674] = 12'b010111110100;
        mem[2675] = 12'b010111110100;
        mem[2676] = 12'b010111110101;
        mem[2677] = 12'b010111110101;
        mem[2678] = 12'b010111110110;
        mem[2679] = 12'b010111110110;
        mem[2680] = 12'b010111110111;
        mem[2681] = 12'b010111110111;
        mem[2682] = 12'b010111110111;
        mem[2683] = 12'b010111111000;
        mem[2684] = 12'b010111111000;
        mem[2685] = 12'b010111111001;
        mem[2686] = 12'b010111111001;
        mem[2687] = 12'b010111111010;
        mem[2688] = 12'b010111111010;
        mem[2689] = 12'b010111111010;
        mem[2690] = 12'b010111111011;
        mem[2691] = 12'b010111111011;
        mem[2692] = 12'b010111111100;
        mem[2693] = 12'b010111111100;
        mem[2694] = 12'b010111111101;
        mem[2695] = 12'b010111111101;
        mem[2696] = 12'b010111111101;
        mem[2697] = 12'b010111111110;
        mem[2698] = 12'b010111111110;
        mem[2699] = 12'b010111111111;
        mem[2700] = 12'b010111111111;
        mem[2701] = 12'b011000000000;
        mem[2702] = 12'b011000000000;
        mem[2703] = 12'b011000000000;
        mem[2704] = 12'b011000000001;
        mem[2705] = 12'b011000000001;
        mem[2706] = 12'b011000000010;
        mem[2707] = 12'b011000000010;
        mem[2708] = 12'b011000000010;
        mem[2709] = 12'b011000000011;
        mem[2710] = 12'b011000000011;
        mem[2711] = 12'b011000000100;
        mem[2712] = 12'b011000000100;
        mem[2713] = 12'b011000000101;
        mem[2714] = 12'b011000000101;
        mem[2715] = 12'b011000000101;
        mem[2716] = 12'b011000000110;
        mem[2717] = 12'b011000000110;
        mem[2718] = 12'b011000000111;
        mem[2719] = 12'b011000000111;
        mem[2720] = 12'b011000001000;
        mem[2721] = 12'b011000001000;
        mem[2722] = 12'b011000001000;
        mem[2723] = 12'b011000001001;
        mem[2724] = 12'b011000001001;
        mem[2725] = 12'b011000001010;
        mem[2726] = 12'b011000001010;
        mem[2727] = 12'b011000001011;
        mem[2728] = 12'b011000001011;
        mem[2729] = 12'b011000001011;
        mem[2730] = 12'b011000001100;
        mem[2731] = 12'b011000001100;
        mem[2732] = 12'b011000001101;
        mem[2733] = 12'b011000001101;
        mem[2734] = 12'b011000001101;
        mem[2735] = 12'b011000001110;
        mem[2736] = 12'b011000001110;
        mem[2737] = 12'b011000001111;
        mem[2738] = 12'b011000001111;
        mem[2739] = 12'b011000010000;
        mem[2740] = 12'b011000010000;
        mem[2741] = 12'b011000010000;
        mem[2742] = 12'b011000010001;
        mem[2743] = 12'b011000010001;
        mem[2744] = 12'b011000010010;
        mem[2745] = 12'b011000010010;
        mem[2746] = 12'b011000010010;
        mem[2747] = 12'b011000010011;
        mem[2748] = 12'b011000010011;
        mem[2749] = 12'b011000010100;
        mem[2750] = 12'b011000010100;
        mem[2751] = 12'b011000010101;
        mem[2752] = 12'b011000010101;
        mem[2753] = 12'b011000010101;
        mem[2754] = 12'b011000010110;
        mem[2755] = 12'b011000010110;
        mem[2756] = 12'b011000010111;
        mem[2757] = 12'b011000010111;
        mem[2758] = 12'b011000011000;
        mem[2759] = 12'b011000011000;
        mem[2760] = 12'b011000011000;
        mem[2761] = 12'b011000011001;
        mem[2762] = 12'b011000011001;
        mem[2763] = 12'b011000011010;
        mem[2764] = 12'b011000011010;
        mem[2765] = 12'b011000011010;
        mem[2766] = 12'b011000011011;
        mem[2767] = 12'b011000011011;
        mem[2768] = 12'b011000011100;
        mem[2769] = 12'b011000011100;
        mem[2770] = 12'b011000011100;
        mem[2771] = 12'b011000011101;
        mem[2772] = 12'b011000011101;
        mem[2773] = 12'b011000011110;
        mem[2774] = 12'b011000011110;
        mem[2775] = 12'b011000011111;
        mem[2776] = 12'b011000011111;
        mem[2777] = 12'b011000011111;
        mem[2778] = 12'b011000100000;
        mem[2779] = 12'b011000100000;
        mem[2780] = 12'b011000100001;
        mem[2781] = 12'b011000100001;
        mem[2782] = 12'b011000100001;
        mem[2783] = 12'b011000100010;
        mem[2784] = 12'b011000100010;
        mem[2785] = 12'b011000100011;
        mem[2786] = 12'b011000100011;
        mem[2787] = 12'b011000100100;
        mem[2788] = 12'b011000100100;
        mem[2789] = 12'b011000100100;
        mem[2790] = 12'b011000100101;
        mem[2791] = 12'b011000100101;
        mem[2792] = 12'b011000100110;
        mem[2793] = 12'b011000100110;
        mem[2794] = 12'b011000100110;
        mem[2795] = 12'b011000100111;
        mem[2796] = 12'b011000100111;
        mem[2797] = 12'b011000101000;
        mem[2798] = 12'b011000101000;
        mem[2799] = 12'b011000101000;
        mem[2800] = 12'b011000101001;
        mem[2801] = 12'b011000101001;
        mem[2802] = 12'b011000101010;
        mem[2803] = 12'b011000101010;
        mem[2804] = 12'b011000101010;
        mem[2805] = 12'b011000101011;
        mem[2806] = 12'b011000101011;
        mem[2807] = 12'b011000101100;
        mem[2808] = 12'b011000101100;
        mem[2809] = 12'b011000101101;
        mem[2810] = 12'b011000101101;
        mem[2811] = 12'b011000101101;
        mem[2812] = 12'b011000101110;
        mem[2813] = 12'b011000101110;
        mem[2814] = 12'b011000101111;
        mem[2815] = 12'b011000101111;
        mem[2816] = 12'b011000101111;
        mem[2817] = 12'b011000110000;
        mem[2818] = 12'b011000110000;
        mem[2819] = 12'b011000110001;
        mem[2820] = 12'b011000110001;
        mem[2821] = 12'b011000110001;
        mem[2822] = 12'b011000110010;
        mem[2823] = 12'b011000110010;
        mem[2824] = 12'b011000110011;
        mem[2825] = 12'b011000110011;
        mem[2826] = 12'b011000110011;
        mem[2827] = 12'b011000110100;
        mem[2828] = 12'b011000110100;
        mem[2829] = 12'b011000110101;
        mem[2830] = 12'b011000110101;
        mem[2831] = 12'b011000110101;
        mem[2832] = 12'b011000110110;
        mem[2833] = 12'b011000110110;
        mem[2834] = 12'b011000110111;
        mem[2835] = 12'b011000110111;
        mem[2836] = 12'b011000111000;
        mem[2837] = 12'b011000111000;
        mem[2838] = 12'b011000111000;
        mem[2839] = 12'b011000111001;
        mem[2840] = 12'b011000111001;
        mem[2841] = 12'b011000111010;
        mem[2842] = 12'b011000111010;
        mem[2843] = 12'b011000111010;
        mem[2844] = 12'b011000111011;
        mem[2845] = 12'b011000111011;
        mem[2846] = 12'b011000111100;
        mem[2847] = 12'b011000111100;
        mem[2848] = 12'b011000111100;
        mem[2849] = 12'b011000111101;
        mem[2850] = 12'b011000111101;
        mem[2851] = 12'b011000111110;
        mem[2852] = 12'b011000111110;
        mem[2853] = 12'b011000111110;
        mem[2854] = 12'b011000111111;
        mem[2855] = 12'b011000111111;
        mem[2856] = 12'b011001000000;
        mem[2857] = 12'b011001000000;
        mem[2858] = 12'b011001000000;
        mem[2859] = 12'b011001000001;
        mem[2860] = 12'b011001000001;
        mem[2861] = 12'b011001000010;
        mem[2862] = 12'b011001000010;
        mem[2863] = 12'b011001000010;
        mem[2864] = 12'b011001000011;
        mem[2865] = 12'b011001000011;
        mem[2866] = 12'b011001000100;
        mem[2867] = 12'b011001000100;
        mem[2868] = 12'b011001000100;
        mem[2869] = 12'b011001000101;
        mem[2870] = 12'b011001000101;
        mem[2871] = 12'b011001000110;
        mem[2872] = 12'b011001000110;
        mem[2873] = 12'b011001000110;
        mem[2874] = 12'b011001000111;
        mem[2875] = 12'b011001000111;
        mem[2876] = 12'b011001001000;
        mem[2877] = 12'b011001001000;
        mem[2878] = 12'b011001001000;
        mem[2879] = 12'b011001001001;
        mem[2880] = 12'b011001001001;
        mem[2881] = 12'b011001001010;
        mem[2882] = 12'b011001001010;
        mem[2883] = 12'b011001001010;
        mem[2884] = 12'b011001001011;
        mem[2885] = 12'b011001001011;
        mem[2886] = 12'b011001001100;
        mem[2887] = 12'b011001001100;
        mem[2888] = 12'b011001001100;
        mem[2889] = 12'b011001001101;
        mem[2890] = 12'b011001001101;
        mem[2891] = 12'b011001001110;
        mem[2892] = 12'b011001001110;
        mem[2893] = 12'b011001001110;
        mem[2894] = 12'b011001001111;
        mem[2895] = 12'b011001001111;
        mem[2896] = 12'b011001001111;
        mem[2897] = 12'b011001010000;
        mem[2898] = 12'b011001010000;
        mem[2899] = 12'b011001010001;
        mem[2900] = 12'b011001010001;
        mem[2901] = 12'b011001010001;
        mem[2902] = 12'b011001010010;
        mem[2903] = 12'b011001010010;
        mem[2904] = 12'b011001010011;
        mem[2905] = 12'b011001010011;
        mem[2906] = 12'b011001010011;
        mem[2907] = 12'b011001010100;
        mem[2908] = 12'b011001010100;
        mem[2909] = 12'b011001010101;
        mem[2910] = 12'b011001010101;
        mem[2911] = 12'b011001010101;
        mem[2912] = 12'b011001010110;
        mem[2913] = 12'b011001010110;
        mem[2914] = 12'b011001010111;
        mem[2915] = 12'b011001010111;
        mem[2916] = 12'b011001010111;
        mem[2917] = 12'b011001011000;
        mem[2918] = 12'b011001011000;
        mem[2919] = 12'b011001011001;
        mem[2920] = 12'b011001011001;
        mem[2921] = 12'b011001011001;
        mem[2922] = 12'b011001011010;
        mem[2923] = 12'b011001011010;
        mem[2924] = 12'b011001011010;
        mem[2925] = 12'b011001011011;
        mem[2926] = 12'b011001011011;
        mem[2927] = 12'b011001011100;
        mem[2928] = 12'b011001011100;
        mem[2929] = 12'b011001011100;
        mem[2930] = 12'b011001011101;
        mem[2931] = 12'b011001011101;
        mem[2932] = 12'b011001011110;
        mem[2933] = 12'b011001011110;
        mem[2934] = 12'b011001011110;
        mem[2935] = 12'b011001011111;
        mem[2936] = 12'b011001011111;
        mem[2937] = 12'b011001100000;
        mem[2938] = 12'b011001100000;
        mem[2939] = 12'b011001100000;
        mem[2940] = 12'b011001100001;
        mem[2941] = 12'b011001100001;
        mem[2942] = 12'b011001100001;
        mem[2943] = 12'b011001100010;
        mem[2944] = 12'b011001100010;
        mem[2945] = 12'b011001100011;
        mem[2946] = 12'b011001100011;
        mem[2947] = 12'b011001100011;
        mem[2948] = 12'b011001100100;
        mem[2949] = 12'b011001100100;
        mem[2950] = 12'b011001100101;
        mem[2951] = 12'b011001100101;
        mem[2952] = 12'b011001100101;
        mem[2953] = 12'b011001100110;
        mem[2954] = 12'b011001100110;
        mem[2955] = 12'b011001100110;
        mem[2956] = 12'b011001100111;
        mem[2957] = 12'b011001100111;
        mem[2958] = 12'b011001101000;
        mem[2959] = 12'b011001101000;
        mem[2960] = 12'b011001101000;
        mem[2961] = 12'b011001101001;
        mem[2962] = 12'b011001101001;
        mem[2963] = 12'b011001101010;
        mem[2964] = 12'b011001101010;
        mem[2965] = 12'b011001101010;
        mem[2966] = 12'b011001101011;
        mem[2967] = 12'b011001101011;
        mem[2968] = 12'b011001101011;
        mem[2969] = 12'b011001101100;
        mem[2970] = 12'b011001101100;
        mem[2971] = 12'b011001101101;
        mem[2972] = 12'b011001101101;
        mem[2973] = 12'b011001101101;
        mem[2974] = 12'b011001101110;
        mem[2975] = 12'b011001101110;
        mem[2976] = 12'b011001101111;
        mem[2977] = 12'b011001101111;
        mem[2978] = 12'b011001101111;
        mem[2979] = 12'b011001110000;
        mem[2980] = 12'b011001110000;
        mem[2981] = 12'b011001110000;
        mem[2982] = 12'b011001110001;
        mem[2983] = 12'b011001110001;
        mem[2984] = 12'b011001110010;
        mem[2985] = 12'b011001110010;
        mem[2986] = 12'b011001110010;
        mem[2987] = 12'b011001110011;
        mem[2988] = 12'b011001110011;
        mem[2989] = 12'b011001110100;
        mem[2990] = 12'b011001110100;
        mem[2991] = 12'b011001110100;
        mem[2992] = 12'b011001110101;
        mem[2993] = 12'b011001110101;
        mem[2994] = 12'b011001110101;
        mem[2995] = 12'b011001110110;
        mem[2996] = 12'b011001110110;
        mem[2997] = 12'b011001110111;
        mem[2998] = 12'b011001110111;
        mem[2999] = 12'b011001110111;
        mem[3000] = 12'b011001111000;
        mem[3001] = 12'b011001111000;
        mem[3002] = 12'b011001111000;
        mem[3003] = 12'b011001111001;
        mem[3004] = 12'b011001111001;
        mem[3005] = 12'b011001111010;
        mem[3006] = 12'b011001111010;
        mem[3007] = 12'b011001111010;
        mem[3008] = 12'b011001111011;
        mem[3009] = 12'b011001111011;
        mem[3010] = 12'b011001111011;
        mem[3011] = 12'b011001111100;
        mem[3012] = 12'b011001111100;
        mem[3013] = 12'b011001111101;
        mem[3014] = 12'b011001111101;
        mem[3015] = 12'b011001111101;
        mem[3016] = 12'b011001111110;
        mem[3017] = 12'b011001111110;
        mem[3018] = 12'b011001111110;
        mem[3019] = 12'b011001111111;
        mem[3020] = 12'b011001111111;
        mem[3021] = 12'b011010000000;
        mem[3022] = 12'b011010000000;
        mem[3023] = 12'b011010000000;
        mem[3024] = 12'b011010000001;
        mem[3025] = 12'b011010000001;
        mem[3026] = 12'b011010000001;
        mem[3027] = 12'b011010000010;
        mem[3028] = 12'b011010000010;
        mem[3029] = 12'b011010000011;
        mem[3030] = 12'b011010000011;
        mem[3031] = 12'b011010000011;
        mem[3032] = 12'b011010000100;
        mem[3033] = 12'b011010000100;
        mem[3034] = 12'b011010000100;
        mem[3035] = 12'b011010000101;
        mem[3036] = 12'b011010000101;
        mem[3037] = 12'b011010000110;
        mem[3038] = 12'b011010000110;
        mem[3039] = 12'b011010000110;
        mem[3040] = 12'b011010000111;
        mem[3041] = 12'b011010000111;
        mem[3042] = 12'b011010000111;
        mem[3043] = 12'b011010001000;
        mem[3044] = 12'b011010001000;
        mem[3045] = 12'b011010001001;
        mem[3046] = 12'b011010001001;
        mem[3047] = 12'b011010001001;
        mem[3048] = 12'b011010001010;
        mem[3049] = 12'b011010001010;
        mem[3050] = 12'b011010001010;
        mem[3051] = 12'b011010001011;
        mem[3052] = 12'b011010001011;
        mem[3053] = 12'b011010001011;
        mem[3054] = 12'b011010001100;
        mem[3055] = 12'b011010001100;
        mem[3056] = 12'b011010001101;
        mem[3057] = 12'b011010001101;
        mem[3058] = 12'b011010001101;
        mem[3059] = 12'b011010001110;
        mem[3060] = 12'b011010001110;
        mem[3061] = 12'b011010001110;
        mem[3062] = 12'b011010001111;
        mem[3063] = 12'b011010001111;
        mem[3064] = 12'b011010010000;
        mem[3065] = 12'b011010010000;
        mem[3066] = 12'b011010010000;
        mem[3067] = 12'b011010010001;
        mem[3068] = 12'b011010010001;
        mem[3069] = 12'b011010010001;
        mem[3070] = 12'b011010010010;
        mem[3071] = 12'b011010010010;
        mem[3072] = 12'b011010010010;
        mem[3073] = 12'b011010010011;
        mem[3074] = 12'b011010010011;
        mem[3075] = 12'b011010010100;
        mem[3076] = 12'b011010010100;
        mem[3077] = 12'b011010010100;
        mem[3078] = 12'b011010010101;
        mem[3079] = 12'b011010010101;
        mem[3080] = 12'b011010010101;
        mem[3081] = 12'b011010010110;
        mem[3082] = 12'b011010010110;
        mem[3083] = 12'b011010010110;
        mem[3084] = 12'b011010010111;
        mem[3085] = 12'b011010010111;
        mem[3086] = 12'b011010011000;
        mem[3087] = 12'b011010011000;
        mem[3088] = 12'b011010011000;
        mem[3089] = 12'b011010011001;
        mem[3090] = 12'b011010011001;
        mem[3091] = 12'b011010011001;
        mem[3092] = 12'b011010011010;
        mem[3093] = 12'b011010011010;
        mem[3094] = 12'b011010011010;
        mem[3095] = 12'b011010011011;
        mem[3096] = 12'b011010011011;
        mem[3097] = 12'b011010011100;
        mem[3098] = 12'b011010011100;
        mem[3099] = 12'b011010011100;
        mem[3100] = 12'b011010011101;
        mem[3101] = 12'b011010011101;
        mem[3102] = 12'b011010011101;
        mem[3103] = 12'b011010011110;
        mem[3104] = 12'b011010011110;
        mem[3105] = 12'b011010011110;
        mem[3106] = 12'b011010011111;
        mem[3107] = 12'b011010011111;
        mem[3108] = 12'b011010100000;
        mem[3109] = 12'b011010100000;
        mem[3110] = 12'b011010100000;
        mem[3111] = 12'b011010100001;
        mem[3112] = 12'b011010100001;
        mem[3113] = 12'b011010100001;
        mem[3114] = 12'b011010100010;
        mem[3115] = 12'b011010100010;
        mem[3116] = 12'b011010100010;
        mem[3117] = 12'b011010100011;
        mem[3118] = 12'b011010100011;
        mem[3119] = 12'b011010100011;
        mem[3120] = 12'b011010100100;
        mem[3121] = 12'b011010100100;
        mem[3122] = 12'b011010100101;
        mem[3123] = 12'b011010100101;
        mem[3124] = 12'b011010100101;
        mem[3125] = 12'b011010100110;
        mem[3126] = 12'b011010100110;
        mem[3127] = 12'b011010100110;
        mem[3128] = 12'b011010100111;
        mem[3129] = 12'b011010100111;
        mem[3130] = 12'b011010100111;
        mem[3131] = 12'b011010101000;
        mem[3132] = 12'b011010101000;
        mem[3133] = 12'b011010101000;
        mem[3134] = 12'b011010101001;
        mem[3135] = 12'b011010101001;
        mem[3136] = 12'b011010101010;
        mem[3137] = 12'b011010101010;
        mem[3138] = 12'b011010101010;
        mem[3139] = 12'b011010101011;
        mem[3140] = 12'b011010101011;
        mem[3141] = 12'b011010101011;
        mem[3142] = 12'b011010101100;
        mem[3143] = 12'b011010101100;
        mem[3144] = 12'b011010101100;
        mem[3145] = 12'b011010101101;
        mem[3146] = 12'b011010101101;
        mem[3147] = 12'b011010101101;
        mem[3148] = 12'b011010101110;
        mem[3149] = 12'b011010101110;
        mem[3150] = 12'b011010101111;
        mem[3151] = 12'b011010101111;
        mem[3152] = 12'b011010101111;
        mem[3153] = 12'b011010110000;
        mem[3154] = 12'b011010110000;
        mem[3155] = 12'b011010110000;
        mem[3156] = 12'b011010110001;
        mem[3157] = 12'b011010110001;
        mem[3158] = 12'b011010110001;
        mem[3159] = 12'b011010110010;
        mem[3160] = 12'b011010110010;
        mem[3161] = 12'b011010110010;
        mem[3162] = 12'b011010110011;
        mem[3163] = 12'b011010110011;
        mem[3164] = 12'b011010110011;
        mem[3165] = 12'b011010110100;
        mem[3166] = 12'b011010110100;
        mem[3167] = 12'b011010110100;
        mem[3168] = 12'b011010110101;
        mem[3169] = 12'b011010110101;
        mem[3170] = 12'b011010110110;
        mem[3171] = 12'b011010110110;
        mem[3172] = 12'b011010110110;
        mem[3173] = 12'b011010110111;
        mem[3174] = 12'b011010110111;
        mem[3175] = 12'b011010110111;
        mem[3176] = 12'b011010111000;
        mem[3177] = 12'b011010111000;
        mem[3178] = 12'b011010111000;
        mem[3179] = 12'b011010111001;
        mem[3180] = 12'b011010111001;
        mem[3181] = 12'b011010111001;
        mem[3182] = 12'b011010111010;
        mem[3183] = 12'b011010111010;
        mem[3184] = 12'b011010111010;
        mem[3185] = 12'b011010111011;
        mem[3186] = 12'b011010111011;
        mem[3187] = 12'b011010111011;
        mem[3188] = 12'b011010111100;
        mem[3189] = 12'b011010111100;
        mem[3190] = 12'b011010111100;
        mem[3191] = 12'b011010111101;
        mem[3192] = 12'b011010111101;
        mem[3193] = 12'b011010111110;
        mem[3194] = 12'b011010111110;
        mem[3195] = 12'b011010111110;
        mem[3196] = 12'b011010111111;
        mem[3197] = 12'b011010111111;
        mem[3198] = 12'b011010111111;
        mem[3199] = 12'b011011000000;
        mem[3200] = 12'b011011000000;
        mem[3201] = 12'b011011000000;
        mem[3202] = 12'b011011000001;
        mem[3203] = 12'b011011000001;
        mem[3204] = 12'b011011000001;
        mem[3205] = 12'b011011000010;
        mem[3206] = 12'b011011000010;
        mem[3207] = 12'b011011000010;
        mem[3208] = 12'b011011000011;
        mem[3209] = 12'b011011000011;
        mem[3210] = 12'b011011000011;
        mem[3211] = 12'b011011000100;
        mem[3212] = 12'b011011000100;
        mem[3213] = 12'b011011000100;
        mem[3214] = 12'b011011000101;
        mem[3215] = 12'b011011000101;
        mem[3216] = 12'b011011000101;
        mem[3217] = 12'b011011000110;
        mem[3218] = 12'b011011000110;
        mem[3219] = 12'b011011000110;
        mem[3220] = 12'b011011000111;
        mem[3221] = 12'b011011000111;
        mem[3222] = 12'b011011000111;
        mem[3223] = 12'b011011001000;
        mem[3224] = 12'b011011001000;
        mem[3225] = 12'b011011001001;
        mem[3226] = 12'b011011001001;
        mem[3227] = 12'b011011001001;
        mem[3228] = 12'b011011001010;
        mem[3229] = 12'b011011001010;
        mem[3230] = 12'b011011001010;
        mem[3231] = 12'b011011001011;
        mem[3232] = 12'b011011001011;
        mem[3233] = 12'b011011001011;
        mem[3234] = 12'b011011001100;
        mem[3235] = 12'b011011001100;
        mem[3236] = 12'b011011001100;
        mem[3237] = 12'b011011001101;
        mem[3238] = 12'b011011001101;
        mem[3239] = 12'b011011001101;
        mem[3240] = 12'b011011001110;
        mem[3241] = 12'b011011001110;
        mem[3242] = 12'b011011001110;
        mem[3243] = 12'b011011001111;
        mem[3244] = 12'b011011001111;
        mem[3245] = 12'b011011001111;
        mem[3246] = 12'b011011010000;
        mem[3247] = 12'b011011010000;
        mem[3248] = 12'b011011010000;
        mem[3249] = 12'b011011010001;
        mem[3250] = 12'b011011010001;
        mem[3251] = 12'b011011010001;
        mem[3252] = 12'b011011010010;
        mem[3253] = 12'b011011010010;
        mem[3254] = 12'b011011010010;
        mem[3255] = 12'b011011010011;
        mem[3256] = 12'b011011010011;
        mem[3257] = 12'b011011010011;
        mem[3258] = 12'b011011010100;
        mem[3259] = 12'b011011010100;
        mem[3260] = 12'b011011010100;
        mem[3261] = 12'b011011010101;
        mem[3262] = 12'b011011010101;
        mem[3263] = 12'b011011010101;
        mem[3264] = 12'b011011010110;
        mem[3265] = 12'b011011010110;
        mem[3266] = 12'b011011010110;
        mem[3267] = 12'b011011010111;
        mem[3268] = 12'b011011010111;
        mem[3269] = 12'b011011010111;
        mem[3270] = 12'b011011011000;
        mem[3271] = 12'b011011011000;
        mem[3272] = 12'b011011011000;
        mem[3273] = 12'b011011011001;
        mem[3274] = 12'b011011011001;
        mem[3275] = 12'b011011011001;
        mem[3276] = 12'b011011011010;
        mem[3277] = 12'b011011011010;
        mem[3278] = 12'b011011011010;
        mem[3279] = 12'b011011011011;
        mem[3280] = 12'b011011011011;
        mem[3281] = 12'b011011011011;
        mem[3282] = 12'b011011011100;
        mem[3283] = 12'b011011011100;
        mem[3284] = 12'b011011011100;
        mem[3285] = 12'b011011011101;
        mem[3286] = 12'b011011011101;
        mem[3287] = 12'b011011011101;
        mem[3288] = 12'b011011011110;
        mem[3289] = 12'b011011011110;
        mem[3290] = 12'b011011011110;
        mem[3291] = 12'b011011011111;
        mem[3292] = 12'b011011011111;
        mem[3293] = 12'b011011011111;
        mem[3294] = 12'b011011100000;
        mem[3295] = 12'b011011100000;
        mem[3296] = 12'b011011100000;
        mem[3297] = 12'b011011100001;
        mem[3298] = 12'b011011100001;
        mem[3299] = 12'b011011100001;
        mem[3300] = 12'b011011100010;
        mem[3301] = 12'b011011100010;
        mem[3302] = 12'b011011100010;
        mem[3303] = 12'b011011100011;
        mem[3304] = 12'b011011100011;
        mem[3305] = 12'b011011100011;
        mem[3306] = 12'b011011100100;
        mem[3307] = 12'b011011100100;
        mem[3308] = 12'b011011100100;
        mem[3309] = 12'b011011100100;
        mem[3310] = 12'b011011100101;
        mem[3311] = 12'b011011100101;
        mem[3312] = 12'b011011100101;
        mem[3313] = 12'b011011100110;
        mem[3314] = 12'b011011100110;
        mem[3315] = 12'b011011100110;
        mem[3316] = 12'b011011100111;
        mem[3317] = 12'b011011100111;
        mem[3318] = 12'b011011100111;
        mem[3319] = 12'b011011101000;
        mem[3320] = 12'b011011101000;
        mem[3321] = 12'b011011101000;
        mem[3322] = 12'b011011101001;
        mem[3323] = 12'b011011101001;
        mem[3324] = 12'b011011101001;
        mem[3325] = 12'b011011101010;
        mem[3326] = 12'b011011101010;
        mem[3327] = 12'b011011101010;
        mem[3328] = 12'b011011101011;
        mem[3329] = 12'b011011101011;
        mem[3330] = 12'b011011101011;
        mem[3331] = 12'b011011101100;
        mem[3332] = 12'b011011101100;
        mem[3333] = 12'b011011101100;
        mem[3334] = 12'b011011101101;
        mem[3335] = 12'b011011101101;
        mem[3336] = 12'b011011101101;
        mem[3337] = 12'b011011101110;
        mem[3338] = 12'b011011101110;
        mem[3339] = 12'b011011101110;
        mem[3340] = 12'b011011101111;
        mem[3341] = 12'b011011101111;
        mem[3342] = 12'b011011101111;
        mem[3343] = 12'b011011101111;
        mem[3344] = 12'b011011110000;
        mem[3345] = 12'b011011110000;
        mem[3346] = 12'b011011110000;
        mem[3347] = 12'b011011110001;
        mem[3348] = 12'b011011110001;
        mem[3349] = 12'b011011110001;
        mem[3350] = 12'b011011110010;
        mem[3351] = 12'b011011110010;
        mem[3352] = 12'b011011110010;
        mem[3353] = 12'b011011110011;
        mem[3354] = 12'b011011110011;
        mem[3355] = 12'b011011110011;
        mem[3356] = 12'b011011110100;
        mem[3357] = 12'b011011110100;
        mem[3358] = 12'b011011110100;
        mem[3359] = 12'b011011110101;
        mem[3360] = 12'b011011110101;
        mem[3361] = 12'b011011110101;
        mem[3362] = 12'b011011110110;
        mem[3363] = 12'b011011110110;
        mem[3364] = 12'b011011110110;
        mem[3365] = 12'b011011110110;
        mem[3366] = 12'b011011110111;
        mem[3367] = 12'b011011110111;
        mem[3368] = 12'b011011110111;
        mem[3369] = 12'b011011111000;
        mem[3370] = 12'b011011111000;
        mem[3371] = 12'b011011111000;
        mem[3372] = 12'b011011111001;
        mem[3373] = 12'b011011111001;
        mem[3374] = 12'b011011111001;
        mem[3375] = 12'b011011111010;
        mem[3376] = 12'b011011111010;
        mem[3377] = 12'b011011111010;
        mem[3378] = 12'b011011111011;
        mem[3379] = 12'b011011111011;
        mem[3380] = 12'b011011111011;
        mem[3381] = 12'b011011111011;
        mem[3382] = 12'b011011111100;
        mem[3383] = 12'b011011111100;
        mem[3384] = 12'b011011111100;
        mem[3385] = 12'b011011111101;
        mem[3386] = 12'b011011111101;
        mem[3387] = 12'b011011111101;
        mem[3388] = 12'b011011111110;
        mem[3389] = 12'b011011111110;
        mem[3390] = 12'b011011111110;
        mem[3391] = 12'b011011111111;
        mem[3392] = 12'b011011111111;
        mem[3393] = 12'b011011111111;
        mem[3394] = 12'b011100000000;
        mem[3395] = 12'b011100000000;
        mem[3396] = 12'b011100000000;
        mem[3397] = 12'b011100000000;
        mem[3398] = 12'b011100000001;
        mem[3399] = 12'b011100000001;
        mem[3400] = 12'b011100000001;
        mem[3401] = 12'b011100000010;
        mem[3402] = 12'b011100000010;
        mem[3403] = 12'b011100000010;
        mem[3404] = 12'b011100000011;
        mem[3405] = 12'b011100000011;
        mem[3406] = 12'b011100000011;
        mem[3407] = 12'b011100000100;
        mem[3408] = 12'b011100000100;
        mem[3409] = 12'b011100000100;
        mem[3410] = 12'b011100000100;
        mem[3411] = 12'b011100000101;
        mem[3412] = 12'b011100000101;
        mem[3413] = 12'b011100000101;
        mem[3414] = 12'b011100000110;
        mem[3415] = 12'b011100000110;
        mem[3416] = 12'b011100000110;
        mem[3417] = 12'b011100000111;
        mem[3418] = 12'b011100000111;
        mem[3419] = 12'b011100000111;
        mem[3420] = 12'b011100001000;
        mem[3421] = 12'b011100001000;
        mem[3422] = 12'b011100001000;
        mem[3423] = 12'b011100001000;
        mem[3424] = 12'b011100001001;
        mem[3425] = 12'b011100001001;
        mem[3426] = 12'b011100001001;
        mem[3427] = 12'b011100001010;
        mem[3428] = 12'b011100001010;
        mem[3429] = 12'b011100001010;
        mem[3430] = 12'b011100001011;
        mem[3431] = 12'b011100001011;
        mem[3432] = 12'b011100001011;
        mem[3433] = 12'b011100001100;
        mem[3434] = 12'b011100001100;
        mem[3435] = 12'b011100001100;
        mem[3436] = 12'b011100001100;
        mem[3437] = 12'b011100001101;
        mem[3438] = 12'b011100001101;
        mem[3439] = 12'b011100001101;
        mem[3440] = 12'b011100001110;
        mem[3441] = 12'b011100001110;
        mem[3442] = 12'b011100001110;
        mem[3443] = 12'b011100001111;
        mem[3444] = 12'b011100001111;
        mem[3445] = 12'b011100001111;
        mem[3446] = 12'b011100001111;
        mem[3447] = 12'b011100010000;
        mem[3448] = 12'b011100010000;
        mem[3449] = 12'b011100010000;
        mem[3450] = 12'b011100010001;
        mem[3451] = 12'b011100010001;
        mem[3452] = 12'b011100010001;
        mem[3453] = 12'b011100010010;
        mem[3454] = 12'b011100010010;
        mem[3455] = 12'b011100010010;
        mem[3456] = 12'b011100010010;
        mem[3457] = 12'b011100010011;
        mem[3458] = 12'b011100010011;
        mem[3459] = 12'b011100010011;
        mem[3460] = 12'b011100010100;
        mem[3461] = 12'b011100010100;
        mem[3462] = 12'b011100010100;
        mem[3463] = 12'b011100010101;
        mem[3464] = 12'b011100010101;
        mem[3465] = 12'b011100010101;
        mem[3466] = 12'b011100010101;
        mem[3467] = 12'b011100010110;
        mem[3468] = 12'b011100010110;
        mem[3469] = 12'b011100010110;
        mem[3470] = 12'b011100010111;
        mem[3471] = 12'b011100010111;
        mem[3472] = 12'b011100010111;
        mem[3473] = 12'b011100011000;
        mem[3474] = 12'b011100011000;
        mem[3475] = 12'b011100011000;
        mem[3476] = 12'b011100011000;
        mem[3477] = 12'b011100011001;
        mem[3478] = 12'b011100011001;
        mem[3479] = 12'b011100011001;
        mem[3480] = 12'b011100011010;
        mem[3481] = 12'b011100011010;
        mem[3482] = 12'b011100011010;
        mem[3483] = 12'b011100011011;
        mem[3484] = 12'b011100011011;
        mem[3485] = 12'b011100011011;
        mem[3486] = 12'b011100011011;
        mem[3487] = 12'b011100011100;
        mem[3488] = 12'b011100011100;
        mem[3489] = 12'b011100011100;
        mem[3490] = 12'b011100011101;
        mem[3491] = 12'b011100011101;
        mem[3492] = 12'b011100011101;
        mem[3493] = 12'b011100011101;
        mem[3494] = 12'b011100011110;
        mem[3495] = 12'b011100011110;
        mem[3496] = 12'b011100011110;
        mem[3497] = 12'b011100011111;
        mem[3498] = 12'b011100011111;
        mem[3499] = 12'b011100011111;
        mem[3500] = 12'b011100011111;
        mem[3501] = 12'b011100100000;
        mem[3502] = 12'b011100100000;
        mem[3503] = 12'b011100100000;
        mem[3504] = 12'b011100100001;
        mem[3505] = 12'b011100100001;
        mem[3506] = 12'b011100100001;
        mem[3507] = 12'b011100100010;
        mem[3508] = 12'b011100100010;
        mem[3509] = 12'b011100100010;
        mem[3510] = 12'b011100100010;
        mem[3511] = 12'b011100100011;
        mem[3512] = 12'b011100100011;
        mem[3513] = 12'b011100100011;
        mem[3514] = 12'b011100100100;
        mem[3515] = 12'b011100100100;
        mem[3516] = 12'b011100100100;
        mem[3517] = 12'b011100100100;
        mem[3518] = 12'b011100100101;
        mem[3519] = 12'b011100100101;
        mem[3520] = 12'b011100100101;
        mem[3521] = 12'b011100100110;
        mem[3522] = 12'b011100100110;
        mem[3523] = 12'b011100100110;
        mem[3524] = 12'b011100100110;
        mem[3525] = 12'b011100100111;
        mem[3526] = 12'b011100100111;
        mem[3527] = 12'b011100100111;
        mem[3528] = 12'b011100101000;
        mem[3529] = 12'b011100101000;
        mem[3530] = 12'b011100101000;
        mem[3531] = 12'b011100101000;
        mem[3532] = 12'b011100101001;
        mem[3533] = 12'b011100101001;
        mem[3534] = 12'b011100101001;
        mem[3535] = 12'b011100101010;
        mem[3536] = 12'b011100101010;
        mem[3537] = 12'b011100101010;
        mem[3538] = 12'b011100101010;
        mem[3539] = 12'b011100101011;
        mem[3540] = 12'b011100101011;
        mem[3541] = 12'b011100101011;
        mem[3542] = 12'b011100101100;
        mem[3543] = 12'b011100101100;
        mem[3544] = 12'b011100101100;
        mem[3545] = 12'b011100101100;
        mem[3546] = 12'b011100101101;
        mem[3547] = 12'b011100101101;
        mem[3548] = 12'b011100101101;
        mem[3549] = 12'b011100101110;
        mem[3550] = 12'b011100101110;
        mem[3551] = 12'b011100101110;
        mem[3552] = 12'b011100101110;
        mem[3553] = 12'b011100101111;
        mem[3554] = 12'b011100101111;
        mem[3555] = 12'b011100101111;
        mem[3556] = 12'b011100110000;
        mem[3557] = 12'b011100110000;
        mem[3558] = 12'b011100110000;
        mem[3559] = 12'b011100110000;
        mem[3560] = 12'b011100110001;
        mem[3561] = 12'b011100110001;
        mem[3562] = 12'b011100110001;
        mem[3563] = 12'b011100110010;
        mem[3564] = 12'b011100110010;
        mem[3565] = 12'b011100110010;
        mem[3566] = 12'b011100110010;
        mem[3567] = 12'b011100110011;
        mem[3568] = 12'b011100110011;
        mem[3569] = 12'b011100110011;
        mem[3570] = 12'b011100110011;
        mem[3571] = 12'b011100110100;
        mem[3572] = 12'b011100110100;
        mem[3573] = 12'b011100110100;
        mem[3574] = 12'b011100110101;
        mem[3575] = 12'b011100110101;
        mem[3576] = 12'b011100110101;
        mem[3577] = 12'b011100110101;
        mem[3578] = 12'b011100110110;
        mem[3579] = 12'b011100110110;
        mem[3580] = 12'b011100110110;
        mem[3581] = 12'b011100110111;
        mem[3582] = 12'b011100110111;
        mem[3583] = 12'b011100110111;
        mem[3584] = 12'b011100110111;
        mem[3585] = 12'b011100111000;
        mem[3586] = 12'b011100111000;
        mem[3587] = 12'b011100111000;
        mem[3588] = 12'b011100111000;
        mem[3589] = 12'b011100111001;
        mem[3590] = 12'b011100111001;
        mem[3591] = 12'b011100111001;
        mem[3592] = 12'b011100111010;
        mem[3593] = 12'b011100111010;
        mem[3594] = 12'b011100111010;
        mem[3595] = 12'b011100111010;
        mem[3596] = 12'b011100111011;
        mem[3597] = 12'b011100111011;
        mem[3598] = 12'b011100111011;
        mem[3599] = 12'b011100111100;
        mem[3600] = 12'b011100111100;
        mem[3601] = 12'b011100111100;
        mem[3602] = 12'b011100111100;
        mem[3603] = 12'b011100111101;
        mem[3604] = 12'b011100111101;
        mem[3605] = 12'b011100111101;
        mem[3606] = 12'b011100111101;
        mem[3607] = 12'b011100111110;
        mem[3608] = 12'b011100111110;
        mem[3609] = 12'b011100111110;
        mem[3610] = 12'b011100111111;
        mem[3611] = 12'b011100111111;
        mem[3612] = 12'b011100111111;
        mem[3613] = 12'b011100111111;
        mem[3614] = 12'b011101000000;
        mem[3615] = 12'b011101000000;
        mem[3616] = 12'b011101000000;
        mem[3617] = 12'b011101000000;
        mem[3618] = 12'b011101000001;
        mem[3619] = 12'b011101000001;
        mem[3620] = 12'b011101000001;
        mem[3621] = 12'b011101000001;
        mem[3622] = 12'b011101000010;
        mem[3623] = 12'b011101000010;
        mem[3624] = 12'b011101000010;
        mem[3625] = 12'b011101000011;
        mem[3626] = 12'b011101000011;
        mem[3627] = 12'b011101000011;
        mem[3628] = 12'b011101000011;
        mem[3629] = 12'b011101000100;
        mem[3630] = 12'b011101000100;
        mem[3631] = 12'b011101000100;
        mem[3632] = 12'b011101000100;
        mem[3633] = 12'b011101000101;
        mem[3634] = 12'b011101000101;
        mem[3635] = 12'b011101000101;
        mem[3636] = 12'b011101000110;
        mem[3637] = 12'b011101000110;
        mem[3638] = 12'b011101000110;
        mem[3639] = 12'b011101000110;
        mem[3640] = 12'b011101000111;
        mem[3641] = 12'b011101000111;
        mem[3642] = 12'b011101000111;
        mem[3643] = 12'b011101000111;
        mem[3644] = 12'b011101001000;
        mem[3645] = 12'b011101001000;
        mem[3646] = 12'b011101001000;
        mem[3647] = 12'b011101001000;
        mem[3648] = 12'b011101001001;
        mem[3649] = 12'b011101001001;
        mem[3650] = 12'b011101001001;
        mem[3651] = 12'b011101001010;
        mem[3652] = 12'b011101001010;
        mem[3653] = 12'b011101001010;
        mem[3654] = 12'b011101001010;
        mem[3655] = 12'b011101001011;
        mem[3656] = 12'b011101001011;
        mem[3657] = 12'b011101001011;
        mem[3658] = 12'b011101001011;
        mem[3659] = 12'b011101001100;
        mem[3660] = 12'b011101001100;
        mem[3661] = 12'b011101001100;
        mem[3662] = 12'b011101001100;
        mem[3663] = 12'b011101001101;
        mem[3664] = 12'b011101001101;
        mem[3665] = 12'b011101001101;
        mem[3666] = 12'b011101001101;
        mem[3667] = 12'b011101001110;
        mem[3668] = 12'b011101001110;
        mem[3669] = 12'b011101001110;
        mem[3670] = 12'b011101001110;
        mem[3671] = 12'b011101001111;
        mem[3672] = 12'b011101001111;
        mem[3673] = 12'b011101001111;
        mem[3674] = 12'b011101010000;
        mem[3675] = 12'b011101010000;
        mem[3676] = 12'b011101010000;
        mem[3677] = 12'b011101010000;
        mem[3678] = 12'b011101010001;
        mem[3679] = 12'b011101010001;
        mem[3680] = 12'b011101010001;
        mem[3681] = 12'b011101010001;
        mem[3682] = 12'b011101010010;
        mem[3683] = 12'b011101010010;
        mem[3684] = 12'b011101010010;
        mem[3685] = 12'b011101010010;
        mem[3686] = 12'b011101010011;
        mem[3687] = 12'b011101010011;
        mem[3688] = 12'b011101010011;
        mem[3689] = 12'b011101010011;
        mem[3690] = 12'b011101010100;
        mem[3691] = 12'b011101010100;
        mem[3692] = 12'b011101010100;
        mem[3693] = 12'b011101010100;
        mem[3694] = 12'b011101010101;
        mem[3695] = 12'b011101010101;
        mem[3696] = 12'b011101010101;
        mem[3697] = 12'b011101010101;
        mem[3698] = 12'b011101010110;
        mem[3699] = 12'b011101010110;
        mem[3700] = 12'b011101010110;
        mem[3701] = 12'b011101010110;
        mem[3702] = 12'b011101010111;
        mem[3703] = 12'b011101010111;
        mem[3704] = 12'b011101010111;
        mem[3705] = 12'b011101011000;
        mem[3706] = 12'b011101011000;
        mem[3707] = 12'b011101011000;
        mem[3708] = 12'b011101011000;
        mem[3709] = 12'b011101011001;
        mem[3710] = 12'b011101011001;
        mem[3711] = 12'b011101011001;
        mem[3712] = 12'b011101011001;
        mem[3713] = 12'b011101011010;
        mem[3714] = 12'b011101011010;
        mem[3715] = 12'b011101011010;
        mem[3716] = 12'b011101011010;
        mem[3717] = 12'b011101011011;
        mem[3718] = 12'b011101011011;
        mem[3719] = 12'b011101011011;
        mem[3720] = 12'b011101011011;
        mem[3721] = 12'b011101011100;
        mem[3722] = 12'b011101011100;
        mem[3723] = 12'b011101011100;
        mem[3724] = 12'b011101011100;
        mem[3725] = 12'b011101011101;
        mem[3726] = 12'b011101011101;
        mem[3727] = 12'b011101011101;
        mem[3728] = 12'b011101011101;
        mem[3729] = 12'b011101011110;
        mem[3730] = 12'b011101011110;
        mem[3731] = 12'b011101011110;
        mem[3732] = 12'b011101011110;
        mem[3733] = 12'b011101011111;
        mem[3734] = 12'b011101011111;
        mem[3735] = 12'b011101011111;
        mem[3736] = 12'b011101011111;
        mem[3737] = 12'b011101100000;
        mem[3738] = 12'b011101100000;
        mem[3739] = 12'b011101100000;
        mem[3740] = 12'b011101100000;
        mem[3741] = 12'b011101100001;
        mem[3742] = 12'b011101100001;
        mem[3743] = 12'b011101100001;
        mem[3744] = 12'b011101100001;
        mem[3745] = 12'b011101100010;
        mem[3746] = 12'b011101100010;
        mem[3747] = 12'b011101100010;
        mem[3748] = 12'b011101100010;
        mem[3749] = 12'b011101100011;
        mem[3750] = 12'b011101100011;
        mem[3751] = 12'b011101100011;
        mem[3752] = 12'b011101100011;
        mem[3753] = 12'b011101100100;
        mem[3754] = 12'b011101100100;
        mem[3755] = 12'b011101100100;
        mem[3756] = 12'b011101100100;
        mem[3757] = 12'b011101100100;
        mem[3758] = 12'b011101100101;
        mem[3759] = 12'b011101100101;
        mem[3760] = 12'b011101100101;
        mem[3761] = 12'b011101100101;
        mem[3762] = 12'b011101100110;
        mem[3763] = 12'b011101100110;
        mem[3764] = 12'b011101100110;
        mem[3765] = 12'b011101100110;
        mem[3766] = 12'b011101100111;
        mem[3767] = 12'b011101100111;
        mem[3768] = 12'b011101100111;
        mem[3769] = 12'b011101100111;
        mem[3770] = 12'b011101101000;
        mem[3771] = 12'b011101101000;
        mem[3772] = 12'b011101101000;
        mem[3773] = 12'b011101101000;
        mem[3774] = 12'b011101101001;
        mem[3775] = 12'b011101101001;
        mem[3776] = 12'b011101101001;
        mem[3777] = 12'b011101101001;
        mem[3778] = 12'b011101101010;
        mem[3779] = 12'b011101101010;
        mem[3780] = 12'b011101101010;
        mem[3781] = 12'b011101101010;
        mem[3782] = 12'b011101101011;
        mem[3783] = 12'b011101101011;
        mem[3784] = 12'b011101101011;
        mem[3785] = 12'b011101101011;
        mem[3786] = 12'b011101101100;
        mem[3787] = 12'b011101101100;
        mem[3788] = 12'b011101101100;
        mem[3789] = 12'b011101101100;
        mem[3790] = 12'b011101101100;
        mem[3791] = 12'b011101101101;
        mem[3792] = 12'b011101101101;
        mem[3793] = 12'b011101101101;
        mem[3794] = 12'b011101101101;
        mem[3795] = 12'b011101101110;
        mem[3796] = 12'b011101101110;
        mem[3797] = 12'b011101101110;
        mem[3798] = 12'b011101101110;
        mem[3799] = 12'b011101101111;
        mem[3800] = 12'b011101101111;
        mem[3801] = 12'b011101101111;
        mem[3802] = 12'b011101101111;
        mem[3803] = 12'b011101110000;
        mem[3804] = 12'b011101110000;
        mem[3805] = 12'b011101110000;
        mem[3806] = 12'b011101110000;
        mem[3807] = 12'b011101110000;
        mem[3808] = 12'b011101110001;
        mem[3809] = 12'b011101110001;
        mem[3810] = 12'b011101110001;
        mem[3811] = 12'b011101110001;
        mem[3812] = 12'b011101110010;
        mem[3813] = 12'b011101110010;
        mem[3814] = 12'b011101110010;
        mem[3815] = 12'b011101110010;
        mem[3816] = 12'b011101110011;
        mem[3817] = 12'b011101110011;
        mem[3818] = 12'b011101110011;
        mem[3819] = 12'b011101110011;
        mem[3820] = 12'b011101110100;
        mem[3821] = 12'b011101110100;
        mem[3822] = 12'b011101110100;
        mem[3823] = 12'b011101110100;
        mem[3824] = 12'b011101110100;
        mem[3825] = 12'b011101110101;
        mem[3826] = 12'b011101110101;
        mem[3827] = 12'b011101110101;
        mem[3828] = 12'b011101110101;
        mem[3829] = 12'b011101110110;
        mem[3830] = 12'b011101110110;
        mem[3831] = 12'b011101110110;
        mem[3832] = 12'b011101110110;
        mem[3833] = 12'b011101110111;
        mem[3834] = 12'b011101110111;
        mem[3835] = 12'b011101110111;
        mem[3836] = 12'b011101110111;
        mem[3837] = 12'b011101110111;
        mem[3838] = 12'b011101111000;
        mem[3839] = 12'b011101111000;
        mem[3840] = 12'b011101111000;
        mem[3841] = 12'b011101111000;
        mem[3842] = 12'b011101111001;
        mem[3843] = 12'b011101111001;
        mem[3844] = 12'b011101111001;
        mem[3845] = 12'b011101111001;
        mem[3846] = 12'b011101111010;
        mem[3847] = 12'b011101111010;
        mem[3848] = 12'b011101111010;
        mem[3849] = 12'b011101111010;
        mem[3850] = 12'b011101111010;
        mem[3851] = 12'b011101111011;
        mem[3852] = 12'b011101111011;
        mem[3853] = 12'b011101111011;
        mem[3854] = 12'b011101111011;
        mem[3855] = 12'b011101111100;
        mem[3856] = 12'b011101111100;
        mem[3857] = 12'b011101111100;
        mem[3858] = 12'b011101111100;
        mem[3859] = 12'b011101111100;
        mem[3860] = 12'b011101111101;
        mem[3861] = 12'b011101111101;
        mem[3862] = 12'b011101111101;
        mem[3863] = 12'b011101111101;
        mem[3864] = 12'b011101111110;
        mem[3865] = 12'b011101111110;
        mem[3866] = 12'b011101111110;
        mem[3867] = 12'b011101111110;
        mem[3868] = 12'b011101111111;
        mem[3869] = 12'b011101111111;
        mem[3870] = 12'b011101111111;
        mem[3871] = 12'b011101111111;
        mem[3872] = 12'b011101111111;
        mem[3873] = 12'b011110000000;
        mem[3874] = 12'b011110000000;
        mem[3875] = 12'b011110000000;
        mem[3876] = 12'b011110000000;
        mem[3877] = 12'b011110000001;
        mem[3878] = 12'b011110000001;
        mem[3879] = 12'b011110000001;
        mem[3880] = 12'b011110000001;
        mem[3881] = 12'b011110000001;
        mem[3882] = 12'b011110000010;
        mem[3883] = 12'b011110000010;
        mem[3884] = 12'b011110000010;
        mem[3885] = 12'b011110000010;
        mem[3886] = 12'b011110000011;
        mem[3887] = 12'b011110000011;
        mem[3888] = 12'b011110000011;
        mem[3889] = 12'b011110000011;
        mem[3890] = 12'b011110000011;
        mem[3891] = 12'b011110000100;
        mem[3892] = 12'b011110000100;
        mem[3893] = 12'b011110000100;
        mem[3894] = 12'b011110000100;
        mem[3895] = 12'b011110000100;
        mem[3896] = 12'b011110000101;
        mem[3897] = 12'b011110000101;
        mem[3898] = 12'b011110000101;
        mem[3899] = 12'b011110000101;
        mem[3900] = 12'b011110000110;
        mem[3901] = 12'b011110000110;
        mem[3902] = 12'b011110000110;
        mem[3903] = 12'b011110000110;
        mem[3904] = 12'b011110000110;
        mem[3905] = 12'b011110000111;
        mem[3906] = 12'b011110000111;
        mem[3907] = 12'b011110000111;
        mem[3908] = 12'b011110000111;
        mem[3909] = 12'b011110001000;
        mem[3910] = 12'b011110001000;
        mem[3911] = 12'b011110001000;
        mem[3912] = 12'b011110001000;
        mem[3913] = 12'b011110001000;
        mem[3914] = 12'b011110001001;
        mem[3915] = 12'b011110001001;
        mem[3916] = 12'b011110001001;
        mem[3917] = 12'b011110001001;
        mem[3918] = 12'b011110001001;
        mem[3919] = 12'b011110001010;
        mem[3920] = 12'b011110001010;
        mem[3921] = 12'b011110001010;
        mem[3922] = 12'b011110001010;
        mem[3923] = 12'b011110001011;
        mem[3924] = 12'b011110001011;
        mem[3925] = 12'b011110001011;
        mem[3926] = 12'b011110001011;
        mem[3927] = 12'b011110001011;
        mem[3928] = 12'b011110001100;
        mem[3929] = 12'b011110001100;
        mem[3930] = 12'b011110001100;
        mem[3931] = 12'b011110001100;
        mem[3932] = 12'b011110001100;
        mem[3933] = 12'b011110001101;
        mem[3934] = 12'b011110001101;
        mem[3935] = 12'b011110001101;
        mem[3936] = 12'b011110001101;
        mem[3937] = 12'b011110001101;
        mem[3938] = 12'b011110001110;
        mem[3939] = 12'b011110001110;
        mem[3940] = 12'b011110001110;
        mem[3941] = 12'b011110001110;
        mem[3942] = 12'b011110001111;
        mem[3943] = 12'b011110001111;
        mem[3944] = 12'b011110001111;
        mem[3945] = 12'b011110001111;
        mem[3946] = 12'b011110001111;
        mem[3947] = 12'b011110010000;
        mem[3948] = 12'b011110010000;
        mem[3949] = 12'b011110010000;
        mem[3950] = 12'b011110010000;
        mem[3951] = 12'b011110010000;
        mem[3952] = 12'b011110010001;
        mem[3953] = 12'b011110010001;
        mem[3954] = 12'b011110010001;
        mem[3955] = 12'b011110010001;
        mem[3956] = 12'b011110010001;
        mem[3957] = 12'b011110010010;
        mem[3958] = 12'b011110010010;
        mem[3959] = 12'b011110010010;
        mem[3960] = 12'b011110010010;
        mem[3961] = 12'b011110010010;
        mem[3962] = 12'b011110010011;
        mem[3963] = 12'b011110010011;
        mem[3964] = 12'b011110010011;
        mem[3965] = 12'b011110010011;
        mem[3966] = 12'b011110010100;
        mem[3967] = 12'b011110010100;
        mem[3968] = 12'b011110010100;
        mem[3969] = 12'b011110010100;
        mem[3970] = 12'b011110010100;
        mem[3971] = 12'b011110010101;
        mem[3972] = 12'b011110010101;
        mem[3973] = 12'b011110010101;
        mem[3974] = 12'b011110010101;
        mem[3975] = 12'b011110010101;
        mem[3976] = 12'b011110010110;
        mem[3977] = 12'b011110010110;
        mem[3978] = 12'b011110010110;
        mem[3979] = 12'b011110010110;
        mem[3980] = 12'b011110010110;
        mem[3981] = 12'b011110010111;
        mem[3982] = 12'b011110010111;
        mem[3983] = 12'b011110010111;
        mem[3984] = 12'b011110010111;
        mem[3985] = 12'b011110010111;
        mem[3986] = 12'b011110011000;
        mem[3987] = 12'b011110011000;
        mem[3988] = 12'b011110011000;
        mem[3989] = 12'b011110011000;
        mem[3990] = 12'b011110011000;
        mem[3991] = 12'b011110011001;
        mem[3992] = 12'b011110011001;
        mem[3993] = 12'b011110011001;
        mem[3994] = 12'b011110011001;
        mem[3995] = 12'b011110011001;
        mem[3996] = 12'b011110011010;
        mem[3997] = 12'b011110011010;
        mem[3998] = 12'b011110011010;
        mem[3999] = 12'b011110011010;
        mem[4000] = 12'b011110011010;
        mem[4001] = 12'b011110011011;
        mem[4002] = 12'b011110011011;
        mem[4003] = 12'b011110011011;
        mem[4004] = 12'b011110011011;
        mem[4005] = 12'b011110011011;
        mem[4006] = 12'b011110011100;
        mem[4007] = 12'b011110011100;
        mem[4008] = 12'b011110011100;
        mem[4009] = 12'b011110011100;
        mem[4010] = 12'b011110011100;
        mem[4011] = 12'b011110011101;
        mem[4012] = 12'b011110011101;
        mem[4013] = 12'b011110011101;
        mem[4014] = 12'b011110011101;
        mem[4015] = 12'b011110011101;
        mem[4016] = 12'b011110011110;
        mem[4017] = 12'b011110011110;
        mem[4018] = 12'b011110011110;
        mem[4019] = 12'b011110011110;
        mem[4020] = 12'b011110011110;
        mem[4021] = 12'b011110011111;
        mem[4022] = 12'b011110011111;
        mem[4023] = 12'b011110011111;
        mem[4024] = 12'b011110011111;
        mem[4025] = 12'b011110011111;
        mem[4026] = 12'b011110011111;
        mem[4027] = 12'b011110100000;
        mem[4028] = 12'b011110100000;
        mem[4029] = 12'b011110100000;
        mem[4030] = 12'b011110100000;
        mem[4031] = 12'b011110100000;
        mem[4032] = 12'b011110100001;
        mem[4033] = 12'b011110100001;
        mem[4034] = 12'b011110100001;
        mem[4035] = 12'b011110100001;
        mem[4036] = 12'b011110100001;
        mem[4037] = 12'b011110100010;
        mem[4038] = 12'b011110100010;
        mem[4039] = 12'b011110100010;
        mem[4040] = 12'b011110100010;
        mem[4041] = 12'b011110100010;
        mem[4042] = 12'b011110100011;
        mem[4043] = 12'b011110100011;
        mem[4044] = 12'b011110100011;
        mem[4045] = 12'b011110100011;
        mem[4046] = 12'b011110100011;
        mem[4047] = 12'b011110100100;
        mem[4048] = 12'b011110100100;
        mem[4049] = 12'b011110100100;
        mem[4050] = 12'b011110100100;
        mem[4051] = 12'b011110100100;
        mem[4052] = 12'b011110100100;
        mem[4053] = 12'b011110100101;
        mem[4054] = 12'b011110100101;
        mem[4055] = 12'b011110100101;
        mem[4056] = 12'b011110100101;
        mem[4057] = 12'b011110100101;
        mem[4058] = 12'b011110100110;
        mem[4059] = 12'b011110100110;
        mem[4060] = 12'b011110100110;
        mem[4061] = 12'b011110100110;
        mem[4062] = 12'b011110100110;
        mem[4063] = 12'b011110100111;
        mem[4064] = 12'b011110100111;
        mem[4065] = 12'b011110100111;
        mem[4066] = 12'b011110100111;
        mem[4067] = 12'b011110100111;
        mem[4068] = 12'b011110100111;
        mem[4069] = 12'b011110101000;
        mem[4070] = 12'b011110101000;
        mem[4071] = 12'b011110101000;
        mem[4072] = 12'b011110101000;
        mem[4073] = 12'b011110101000;
        mem[4074] = 12'b011110101001;
        mem[4075] = 12'b011110101001;
        mem[4076] = 12'b011110101001;
        mem[4077] = 12'b011110101001;
        mem[4078] = 12'b011110101001;
        mem[4079] = 12'b011110101001;
        mem[4080] = 12'b011110101010;
        mem[4081] = 12'b011110101010;
        mem[4082] = 12'b011110101010;
        mem[4083] = 12'b011110101010;
        mem[4084] = 12'b011110101010;
        mem[4085] = 12'b011110101011;
        mem[4086] = 12'b011110101011;
        mem[4087] = 12'b011110101011;
        mem[4088] = 12'b011110101011;
        mem[4089] = 12'b011110101011;
        mem[4090] = 12'b011110101011;
        mem[4091] = 12'b011110101100;
        mem[4092] = 12'b011110101100;
        mem[4093] = 12'b011110101100;
        mem[4094] = 12'b011110101100;
        mem[4095] = 12'b011110101100;
        mem[4096] = 12'b011110101101;
        mem[4097] = 12'b011110101101;
        mem[4098] = 12'b011110101101;
        mem[4099] = 12'b011110101101;
        mem[4100] = 12'b011110101101;
        mem[4101] = 12'b011110101101;
        mem[4102] = 12'b011110101110;
        mem[4103] = 12'b011110101110;
        mem[4104] = 12'b011110101110;
        mem[4105] = 12'b011110101110;
        mem[4106] = 12'b011110101110;
        mem[4107] = 12'b011110101111;
        mem[4108] = 12'b011110101111;
        mem[4109] = 12'b011110101111;
        mem[4110] = 12'b011110101111;
        mem[4111] = 12'b011110101111;
        mem[4112] = 12'b011110101111;
        mem[4113] = 12'b011110110000;
        mem[4114] = 12'b011110110000;
        mem[4115] = 12'b011110110000;
        mem[4116] = 12'b011110110000;
        mem[4117] = 12'b011110110000;
        mem[4118] = 12'b011110110000;
        mem[4119] = 12'b011110110001;
        mem[4120] = 12'b011110110001;
        mem[4121] = 12'b011110110001;
        mem[4122] = 12'b011110110001;
        mem[4123] = 12'b011110110001;
        mem[4124] = 12'b011110110010;
        mem[4125] = 12'b011110110010;
        mem[4126] = 12'b011110110010;
        mem[4127] = 12'b011110110010;
        mem[4128] = 12'b011110110010;
        mem[4129] = 12'b011110110010;
        mem[4130] = 12'b011110110011;
        mem[4131] = 12'b011110110011;
        mem[4132] = 12'b011110110011;
        mem[4133] = 12'b011110110011;
        mem[4134] = 12'b011110110011;
        mem[4135] = 12'b011110110011;
        mem[4136] = 12'b011110110100;
        mem[4137] = 12'b011110110100;
        mem[4138] = 12'b011110110100;
        mem[4139] = 12'b011110110100;
        mem[4140] = 12'b011110110100;
        mem[4141] = 12'b011110110100;
        mem[4142] = 12'b011110110101;
        mem[4143] = 12'b011110110101;
        mem[4144] = 12'b011110110101;
        mem[4145] = 12'b011110110101;
        mem[4146] = 12'b011110110101;
        mem[4147] = 12'b011110110110;
        mem[4148] = 12'b011110110110;
        mem[4149] = 12'b011110110110;
        mem[4150] = 12'b011110110110;
        mem[4151] = 12'b011110110110;
        mem[4152] = 12'b011110110110;
        mem[4153] = 12'b011110110111;
        mem[4154] = 12'b011110110111;
        mem[4155] = 12'b011110110111;
        mem[4156] = 12'b011110110111;
        mem[4157] = 12'b011110110111;
        mem[4158] = 12'b011110110111;
        mem[4159] = 12'b011110111000;
        mem[4160] = 12'b011110111000;
        mem[4161] = 12'b011110111000;
        mem[4162] = 12'b011110111000;
        mem[4163] = 12'b011110111000;
        mem[4164] = 12'b011110111000;
        mem[4165] = 12'b011110111001;
        mem[4166] = 12'b011110111001;
        mem[4167] = 12'b011110111001;
        mem[4168] = 12'b011110111001;
        mem[4169] = 12'b011110111001;
        mem[4170] = 12'b011110111001;
        mem[4171] = 12'b011110111010;
        mem[4172] = 12'b011110111010;
        mem[4173] = 12'b011110111010;
        mem[4174] = 12'b011110111010;
        mem[4175] = 12'b011110111010;
        mem[4176] = 12'b011110111010;
        mem[4177] = 12'b011110111011;
        mem[4178] = 12'b011110111011;
        mem[4179] = 12'b011110111011;
        mem[4180] = 12'b011110111011;
        mem[4181] = 12'b011110111011;
        mem[4182] = 12'b011110111011;
        mem[4183] = 12'b011110111100;
        mem[4184] = 12'b011110111100;
        mem[4185] = 12'b011110111100;
        mem[4186] = 12'b011110111100;
        mem[4187] = 12'b011110111100;
        mem[4188] = 12'b011110111100;
        mem[4189] = 12'b011110111100;
        mem[4190] = 12'b011110111101;
        mem[4191] = 12'b011110111101;
        mem[4192] = 12'b011110111101;
        mem[4193] = 12'b011110111101;
        mem[4194] = 12'b011110111101;
        mem[4195] = 12'b011110111101;
        mem[4196] = 12'b011110111110;
        mem[4197] = 12'b011110111110;
        mem[4198] = 12'b011110111110;
        mem[4199] = 12'b011110111110;
        mem[4200] = 12'b011110111110;
        mem[4201] = 12'b011110111110;
        mem[4202] = 12'b011110111111;
        mem[4203] = 12'b011110111111;
        mem[4204] = 12'b011110111111;
        mem[4205] = 12'b011110111111;
        mem[4206] = 12'b011110111111;
        mem[4207] = 12'b011110111111;
        mem[4208] = 12'b011111000000;
        mem[4209] = 12'b011111000000;
        mem[4210] = 12'b011111000000;
        mem[4211] = 12'b011111000000;
        mem[4212] = 12'b011111000000;
        mem[4213] = 12'b011111000000;
        mem[4214] = 12'b011111000000;
        mem[4215] = 12'b011111000001;
        mem[4216] = 12'b011111000001;
        mem[4217] = 12'b011111000001;
        mem[4218] = 12'b011111000001;
        mem[4219] = 12'b011111000001;
        mem[4220] = 12'b011111000001;
        mem[4221] = 12'b011111000010;
        mem[4222] = 12'b011111000010;
        mem[4223] = 12'b011111000010;
        mem[4224] = 12'b011111000010;
        mem[4225] = 12'b011111000010;
        mem[4226] = 12'b011111000010;
        mem[4227] = 12'b011111000011;
        mem[4228] = 12'b011111000011;
        mem[4229] = 12'b011111000011;
        mem[4230] = 12'b011111000011;
        mem[4231] = 12'b011111000011;
        mem[4232] = 12'b011111000011;
        mem[4233] = 12'b011111000011;
        mem[4234] = 12'b011111000100;
        mem[4235] = 12'b011111000100;
        mem[4236] = 12'b011111000100;
        mem[4237] = 12'b011111000100;
        mem[4238] = 12'b011111000100;
        mem[4239] = 12'b011111000100;
        mem[4240] = 12'b011111000100;
        mem[4241] = 12'b011111000101;
        mem[4242] = 12'b011111000101;
        mem[4243] = 12'b011111000101;
        mem[4244] = 12'b011111000101;
        mem[4245] = 12'b011111000101;
        mem[4246] = 12'b011111000101;
        mem[4247] = 12'b011111000110;
        mem[4248] = 12'b011111000110;
        mem[4249] = 12'b011111000110;
        mem[4250] = 12'b011111000110;
        mem[4251] = 12'b011111000110;
        mem[4252] = 12'b011111000110;
        mem[4253] = 12'b011111000110;
        mem[4254] = 12'b011111000111;
        mem[4255] = 12'b011111000111;
        mem[4256] = 12'b011111000111;
        mem[4257] = 12'b011111000111;
        mem[4258] = 12'b011111000111;
        mem[4259] = 12'b011111000111;
        mem[4260] = 12'b011111000111;
        mem[4261] = 12'b011111001000;
        mem[4262] = 12'b011111001000;
        mem[4263] = 12'b011111001000;
        mem[4264] = 12'b011111001000;
        mem[4265] = 12'b011111001000;
        mem[4266] = 12'b011111001000;
        mem[4267] = 12'b011111001001;
        mem[4268] = 12'b011111001001;
        mem[4269] = 12'b011111001001;
        mem[4270] = 12'b011111001001;
        mem[4271] = 12'b011111001001;
        mem[4272] = 12'b011111001001;
        mem[4273] = 12'b011111001001;
        mem[4274] = 12'b011111001010;
        mem[4275] = 12'b011111001010;
        mem[4276] = 12'b011111001010;
        mem[4277] = 12'b011111001010;
        mem[4278] = 12'b011111001010;
        mem[4279] = 12'b011111001010;
        mem[4280] = 12'b011111001010;
        mem[4281] = 12'b011111001011;
        mem[4282] = 12'b011111001011;
        mem[4283] = 12'b011111001011;
        mem[4284] = 12'b011111001011;
        mem[4285] = 12'b011111001011;
        mem[4286] = 12'b011111001011;
        mem[4287] = 12'b011111001011;
        mem[4288] = 12'b011111001100;
        mem[4289] = 12'b011111001100;
        mem[4290] = 12'b011111001100;
        mem[4291] = 12'b011111001100;
        mem[4292] = 12'b011111001100;
        mem[4293] = 12'b011111001100;
        mem[4294] = 12'b011111001100;
        mem[4295] = 12'b011111001101;
        mem[4296] = 12'b011111001101;
        mem[4297] = 12'b011111001101;
        mem[4298] = 12'b011111001101;
        mem[4299] = 12'b011111001101;
        mem[4300] = 12'b011111001101;
        mem[4301] = 12'b011111001101;
        mem[4302] = 12'b011111001110;
        mem[4303] = 12'b011111001110;
        mem[4304] = 12'b011111001110;
        mem[4305] = 12'b011111001110;
        mem[4306] = 12'b011111001110;
        mem[4307] = 12'b011111001110;
        mem[4308] = 12'b011111001110;
        mem[4309] = 12'b011111001111;
        mem[4310] = 12'b011111001111;
        mem[4311] = 12'b011111001111;
        mem[4312] = 12'b011111001111;
        mem[4313] = 12'b011111001111;
        mem[4314] = 12'b011111001111;
        mem[4315] = 12'b011111001111;
        mem[4316] = 12'b011111001111;
        mem[4317] = 12'b011111010000;
        mem[4318] = 12'b011111010000;
        mem[4319] = 12'b011111010000;
        mem[4320] = 12'b011111010000;
        mem[4321] = 12'b011111010000;
        mem[4322] = 12'b011111010000;
        mem[4323] = 12'b011111010000;
        mem[4324] = 12'b011111010001;
        mem[4325] = 12'b011111010001;
        mem[4326] = 12'b011111010001;
        mem[4327] = 12'b011111010001;
        mem[4328] = 12'b011111010001;
        mem[4329] = 12'b011111010001;
        mem[4330] = 12'b011111010001;
        mem[4331] = 12'b011111010010;
        mem[4332] = 12'b011111010010;
        mem[4333] = 12'b011111010010;
        mem[4334] = 12'b011111010010;
        mem[4335] = 12'b011111010010;
        mem[4336] = 12'b011111010010;
        mem[4337] = 12'b011111010010;
        mem[4338] = 12'b011111010010;
        mem[4339] = 12'b011111010011;
        mem[4340] = 12'b011111010011;
        mem[4341] = 12'b011111010011;
        mem[4342] = 12'b011111010011;
        mem[4343] = 12'b011111010011;
        mem[4344] = 12'b011111010011;
        mem[4345] = 12'b011111010011;
        mem[4346] = 12'b011111010100;
        mem[4347] = 12'b011111010100;
        mem[4348] = 12'b011111010100;
        mem[4349] = 12'b011111010100;
        mem[4350] = 12'b011111010100;
        mem[4351] = 12'b011111010100;
        mem[4352] = 12'b011111010100;
        mem[4353] = 12'b011111010100;
        mem[4354] = 12'b011111010101;
        mem[4355] = 12'b011111010101;
        mem[4356] = 12'b011111010101;
        mem[4357] = 12'b011111010101;
        mem[4358] = 12'b011111010101;
        mem[4359] = 12'b011111010101;
        mem[4360] = 12'b011111010101;
        mem[4361] = 12'b011111010101;
        mem[4362] = 12'b011111010110;
        mem[4363] = 12'b011111010110;
        mem[4364] = 12'b011111010110;
        mem[4365] = 12'b011111010110;
        mem[4366] = 12'b011111010110;
        mem[4367] = 12'b011111010110;
        mem[4368] = 12'b011111010110;
        mem[4369] = 12'b011111010110;
        mem[4370] = 12'b011111010111;
        mem[4371] = 12'b011111010111;
        mem[4372] = 12'b011111010111;
        mem[4373] = 12'b011111010111;
        mem[4374] = 12'b011111010111;
        mem[4375] = 12'b011111010111;
        mem[4376] = 12'b011111010111;
        mem[4377] = 12'b011111010111;
        mem[4378] = 12'b011111011000;
        mem[4379] = 12'b011111011000;
        mem[4380] = 12'b011111011000;
        mem[4381] = 12'b011111011000;
        mem[4382] = 12'b011111011000;
        mem[4383] = 12'b011111011000;
        mem[4384] = 12'b011111011000;
        mem[4385] = 12'b011111011000;
        mem[4386] = 12'b011111011001;
        mem[4387] = 12'b011111011001;
        mem[4388] = 12'b011111011001;
        mem[4389] = 12'b011111011001;
        mem[4390] = 12'b011111011001;
        mem[4391] = 12'b011111011001;
        mem[4392] = 12'b011111011001;
        mem[4393] = 12'b011111011001;
        mem[4394] = 12'b011111011010;
        mem[4395] = 12'b011111011010;
        mem[4396] = 12'b011111011010;
        mem[4397] = 12'b011111011010;
        mem[4398] = 12'b011111011010;
        mem[4399] = 12'b011111011010;
        mem[4400] = 12'b011111011010;
        mem[4401] = 12'b011111011010;
        mem[4402] = 12'b011111011011;
        mem[4403] = 12'b011111011011;
        mem[4404] = 12'b011111011011;
        mem[4405] = 12'b011111011011;
        mem[4406] = 12'b011111011011;
        mem[4407] = 12'b011111011011;
        mem[4408] = 12'b011111011011;
        mem[4409] = 12'b011111011011;
        mem[4410] = 12'b011111011011;
        mem[4411] = 12'b011111011100;
        mem[4412] = 12'b011111011100;
        mem[4413] = 12'b011111011100;
        mem[4414] = 12'b011111011100;
        mem[4415] = 12'b011111011100;
        mem[4416] = 12'b011111011100;
        mem[4417] = 12'b011111011100;
        mem[4418] = 12'b011111011100;
        mem[4419] = 12'b011111011101;
        mem[4420] = 12'b011111011101;
        mem[4421] = 12'b011111011101;
        mem[4422] = 12'b011111011101;
        mem[4423] = 12'b011111011101;
        mem[4424] = 12'b011111011101;
        mem[4425] = 12'b011111011101;
        mem[4426] = 12'b011111011101;
        mem[4427] = 12'b011111011101;
        mem[4428] = 12'b011111011110;
        mem[4429] = 12'b011111011110;
        mem[4430] = 12'b011111011110;
        mem[4431] = 12'b011111011110;
        mem[4432] = 12'b011111011110;
        mem[4433] = 12'b011111011110;
        mem[4434] = 12'b011111011110;
        mem[4435] = 12'b011111011110;
        mem[4436] = 12'b011111011111;
        mem[4437] = 12'b011111011111;
        mem[4438] = 12'b011111011111;
        mem[4439] = 12'b011111011111;
        mem[4440] = 12'b011111011111;
        mem[4441] = 12'b011111011111;
        mem[4442] = 12'b011111011111;
        mem[4443] = 12'b011111011111;
        mem[4444] = 12'b011111011111;
        mem[4445] = 12'b011111100000;
        mem[4446] = 12'b011111100000;
        mem[4447] = 12'b011111100000;
        mem[4448] = 12'b011111100000;
        mem[4449] = 12'b011111100000;
        mem[4450] = 12'b011111100000;
        mem[4451] = 12'b011111100000;
        mem[4452] = 12'b011111100000;
        mem[4453] = 12'b011111100000;
        mem[4454] = 12'b011111100001;
        mem[4455] = 12'b011111100001;
        mem[4456] = 12'b011111100001;
        mem[4457] = 12'b011111100001;
        mem[4458] = 12'b011111100001;
        mem[4459] = 12'b011111100001;
        mem[4460] = 12'b011111100001;
        mem[4461] = 12'b011111100001;
        mem[4462] = 12'b011111100001;
        mem[4463] = 12'b011111100001;
        mem[4464] = 12'b011111100010;
        mem[4465] = 12'b011111100010;
        mem[4466] = 12'b011111100010;
        mem[4467] = 12'b011111100010;
        mem[4468] = 12'b011111100010;
        mem[4469] = 12'b011111100010;
        mem[4470] = 12'b011111100010;
        mem[4471] = 12'b011111100010;
        mem[4472] = 12'b011111100010;
        mem[4473] = 12'b011111100011;
        mem[4474] = 12'b011111100011;
        mem[4475] = 12'b011111100011;
        mem[4476] = 12'b011111100011;
        mem[4477] = 12'b011111100011;
        mem[4478] = 12'b011111100011;
        mem[4479] = 12'b011111100011;
        mem[4480] = 12'b011111100011;
        mem[4481] = 12'b011111100011;
        mem[4482] = 12'b011111100100;
        mem[4483] = 12'b011111100100;
        mem[4484] = 12'b011111100100;
        mem[4485] = 12'b011111100100;
        mem[4486] = 12'b011111100100;
        mem[4487] = 12'b011111100100;
        mem[4488] = 12'b011111100100;
        mem[4489] = 12'b011111100100;
        mem[4490] = 12'b011111100100;
        mem[4491] = 12'b011111100100;
        mem[4492] = 12'b011111100101;
        mem[4493] = 12'b011111100101;
        mem[4494] = 12'b011111100101;
        mem[4495] = 12'b011111100101;
        mem[4496] = 12'b011111100101;
        mem[4497] = 12'b011111100101;
        mem[4498] = 12'b011111100101;
        mem[4499] = 12'b011111100101;
        mem[4500] = 12'b011111100101;
        mem[4501] = 12'b011111100101;
        mem[4502] = 12'b011111100110;
        mem[4503] = 12'b011111100110;
        mem[4504] = 12'b011111100110;
        mem[4505] = 12'b011111100110;
        mem[4506] = 12'b011111100110;
        mem[4507] = 12'b011111100110;
        mem[4508] = 12'b011111100110;
        mem[4509] = 12'b011111100110;
        mem[4510] = 12'b011111100110;
        mem[4511] = 12'b011111100110;
        mem[4512] = 12'b011111100111;
        mem[4513] = 12'b011111100111;
        mem[4514] = 12'b011111100111;
        mem[4515] = 12'b011111100111;
        mem[4516] = 12'b011111100111;
        mem[4517] = 12'b011111100111;
        mem[4518] = 12'b011111100111;
        mem[4519] = 12'b011111100111;
        mem[4520] = 12'b011111100111;
        mem[4521] = 12'b011111100111;
        mem[4522] = 12'b011111101000;
        mem[4523] = 12'b011111101000;
        mem[4524] = 12'b011111101000;
        mem[4525] = 12'b011111101000;
        mem[4526] = 12'b011111101000;
        mem[4527] = 12'b011111101000;
        mem[4528] = 12'b011111101000;
        mem[4529] = 12'b011111101000;
        mem[4530] = 12'b011111101000;
        mem[4531] = 12'b011111101000;
        mem[4532] = 12'b011111101000;
        mem[4533] = 12'b011111101001;
        mem[4534] = 12'b011111101001;
        mem[4535] = 12'b011111101001;
        mem[4536] = 12'b011111101001;
        mem[4537] = 12'b011111101001;
        mem[4538] = 12'b011111101001;
        mem[4539] = 12'b011111101001;
        mem[4540] = 12'b011111101001;
        mem[4541] = 12'b011111101001;
        mem[4542] = 12'b011111101001;
        mem[4543] = 12'b011111101001;
        mem[4544] = 12'b011111101010;
        mem[4545] = 12'b011111101010;
        mem[4546] = 12'b011111101010;
        mem[4547] = 12'b011111101010;
        mem[4548] = 12'b011111101010;
        mem[4549] = 12'b011111101010;
        mem[4550] = 12'b011111101010;
        mem[4551] = 12'b011111101010;
        mem[4552] = 12'b011111101010;
        mem[4553] = 12'b011111101010;
        mem[4554] = 12'b011111101010;
        mem[4555] = 12'b011111101011;
        mem[4556] = 12'b011111101011;
        mem[4557] = 12'b011111101011;
        mem[4558] = 12'b011111101011;
        mem[4559] = 12'b011111101011;
        mem[4560] = 12'b011111101011;
        mem[4561] = 12'b011111101011;
        mem[4562] = 12'b011111101011;
        mem[4563] = 12'b011111101011;
        mem[4564] = 12'b011111101011;
        mem[4565] = 12'b011111101011;
        mem[4566] = 12'b011111101100;
        mem[4567] = 12'b011111101100;
        mem[4568] = 12'b011111101100;
        mem[4569] = 12'b011111101100;
        mem[4570] = 12'b011111101100;
        mem[4571] = 12'b011111101100;
        mem[4572] = 12'b011111101100;
        mem[4573] = 12'b011111101100;
        mem[4574] = 12'b011111101100;
        mem[4575] = 12'b011111101100;
        mem[4576] = 12'b011111101100;
        mem[4577] = 12'b011111101100;
        mem[4578] = 12'b011111101101;
        mem[4579] = 12'b011111101101;
        mem[4580] = 12'b011111101101;
        mem[4581] = 12'b011111101101;
        mem[4582] = 12'b011111101101;
        mem[4583] = 12'b011111101101;
        mem[4584] = 12'b011111101101;
        mem[4585] = 12'b011111101101;
        mem[4586] = 12'b011111101101;
        mem[4587] = 12'b011111101101;
        mem[4588] = 12'b011111101101;
        mem[4589] = 12'b011111101101;
        mem[4590] = 12'b011111101110;
        mem[4591] = 12'b011111101110;
        mem[4592] = 12'b011111101110;
        mem[4593] = 12'b011111101110;
        mem[4594] = 12'b011111101110;
        mem[4595] = 12'b011111101110;
        mem[4596] = 12'b011111101110;
        mem[4597] = 12'b011111101110;
        mem[4598] = 12'b011111101110;
        mem[4599] = 12'b011111101110;
        mem[4600] = 12'b011111101110;
        mem[4601] = 12'b011111101110;
        mem[4602] = 12'b011111101111;
        mem[4603] = 12'b011111101111;
        mem[4604] = 12'b011111101111;
        mem[4605] = 12'b011111101111;
        mem[4606] = 12'b011111101111;
        mem[4607] = 12'b011111101111;
        mem[4608] = 12'b011111101111;
        mem[4609] = 12'b011111101111;
        mem[4610] = 12'b011111101111;
        mem[4611] = 12'b011111101111;
        mem[4612] = 12'b011111101111;
        mem[4613] = 12'b011111101111;
        mem[4614] = 12'b011111110000;
        mem[4615] = 12'b011111110000;
        mem[4616] = 12'b011111110000;
        mem[4617] = 12'b011111110000;
        mem[4618] = 12'b011111110000;
        mem[4619] = 12'b011111110000;
        mem[4620] = 12'b011111110000;
        mem[4621] = 12'b011111110000;
        mem[4622] = 12'b011111110000;
        mem[4623] = 12'b011111110000;
        mem[4624] = 12'b011111110000;
        mem[4625] = 12'b011111110000;
        mem[4626] = 12'b011111110000;
        mem[4627] = 12'b011111110000;
        mem[4628] = 12'b011111110001;
        mem[4629] = 12'b011111110001;
        mem[4630] = 12'b011111110001;
        mem[4631] = 12'b011111110001;
        mem[4632] = 12'b011111110001;
        mem[4633] = 12'b011111110001;
        mem[4634] = 12'b011111110001;
        mem[4635] = 12'b011111110001;
        mem[4636] = 12'b011111110001;
        mem[4637] = 12'b011111110001;
        mem[4638] = 12'b011111110001;
        mem[4639] = 12'b011111110001;
        mem[4640] = 12'b011111110001;
        mem[4641] = 12'b011111110010;
        mem[4642] = 12'b011111110010;
        mem[4643] = 12'b011111110010;
        mem[4644] = 12'b011111110010;
        mem[4645] = 12'b011111110010;
        mem[4646] = 12'b011111110010;
        mem[4647] = 12'b011111110010;
        mem[4648] = 12'b011111110010;
        mem[4649] = 12'b011111110010;
        mem[4650] = 12'b011111110010;
        mem[4651] = 12'b011111110010;
        mem[4652] = 12'b011111110010;
        mem[4653] = 12'b011111110010;
        mem[4654] = 12'b011111110010;
        mem[4655] = 12'b011111110011;
        mem[4656] = 12'b011111110011;
        mem[4657] = 12'b011111110011;
        mem[4658] = 12'b011111110011;
        mem[4659] = 12'b011111110011;
        mem[4660] = 12'b011111110011;
        mem[4661] = 12'b011111110011;
        mem[4662] = 12'b011111110011;
        mem[4663] = 12'b011111110011;
        mem[4664] = 12'b011111110011;
        mem[4665] = 12'b011111110011;
        mem[4666] = 12'b011111110011;
        mem[4667] = 12'b011111110011;
        mem[4668] = 12'b011111110011;
        mem[4669] = 12'b011111110011;
        mem[4670] = 12'b011111110100;
        mem[4671] = 12'b011111110100;
        mem[4672] = 12'b011111110100;
        mem[4673] = 12'b011111110100;
        mem[4674] = 12'b011111110100;
        mem[4675] = 12'b011111110100;
        mem[4676] = 12'b011111110100;
        mem[4677] = 12'b011111110100;
        mem[4678] = 12'b011111110100;
        mem[4679] = 12'b011111110100;
        mem[4680] = 12'b011111110100;
        mem[4681] = 12'b011111110100;
        mem[4682] = 12'b011111110100;
        mem[4683] = 12'b011111110100;
        mem[4684] = 12'b011111110100;
        mem[4685] = 12'b011111110101;
        mem[4686] = 12'b011111110101;
        mem[4687] = 12'b011111110101;
        mem[4688] = 12'b011111110101;
        mem[4689] = 12'b011111110101;
        mem[4690] = 12'b011111110101;
        mem[4691] = 12'b011111110101;
        mem[4692] = 12'b011111110101;
        mem[4693] = 12'b011111110101;
        mem[4694] = 12'b011111110101;
        mem[4695] = 12'b011111110101;
        mem[4696] = 12'b011111110101;
        mem[4697] = 12'b011111110101;
        mem[4698] = 12'b011111110101;
        mem[4699] = 12'b011111110101;
        mem[4700] = 12'b011111110101;
        mem[4701] = 12'b011111110110;
        mem[4702] = 12'b011111110110;
        mem[4703] = 12'b011111110110;
        mem[4704] = 12'b011111110110;
        mem[4705] = 12'b011111110110;
        mem[4706] = 12'b011111110110;
        mem[4707] = 12'b011111110110;
        mem[4708] = 12'b011111110110;
        mem[4709] = 12'b011111110110;
        mem[4710] = 12'b011111110110;
        mem[4711] = 12'b011111110110;
        mem[4712] = 12'b011111110110;
        mem[4713] = 12'b011111110110;
        mem[4714] = 12'b011111110110;
        mem[4715] = 12'b011111110110;
        mem[4716] = 12'b011111110110;
        mem[4717] = 12'b011111110110;
        mem[4718] = 12'b011111110110;
        mem[4719] = 12'b011111110111;
        mem[4720] = 12'b011111110111;
        mem[4721] = 12'b011111110111;
        mem[4722] = 12'b011111110111;
        mem[4723] = 12'b011111110111;
        mem[4724] = 12'b011111110111;
        mem[4725] = 12'b011111110111;
        mem[4726] = 12'b011111110111;
        mem[4727] = 12'b011111110111;
        mem[4728] = 12'b011111110111;
        mem[4729] = 12'b011111110111;
        mem[4730] = 12'b011111110111;
        mem[4731] = 12'b011111110111;
        mem[4732] = 12'b011111110111;
        mem[4733] = 12'b011111110111;
        mem[4734] = 12'b011111110111;
        mem[4735] = 12'b011111110111;
        mem[4736] = 12'b011111110111;
        mem[4737] = 12'b011111111000;
        mem[4738] = 12'b011111111000;
        mem[4739] = 12'b011111111000;
        mem[4740] = 12'b011111111000;
        mem[4741] = 12'b011111111000;
        mem[4742] = 12'b011111111000;
        mem[4743] = 12'b011111111000;
        mem[4744] = 12'b011111111000;
        mem[4745] = 12'b011111111000;
        mem[4746] = 12'b011111111000;
        mem[4747] = 12'b011111111000;
        mem[4748] = 12'b011111111000;
        mem[4749] = 12'b011111111000;
        mem[4750] = 12'b011111111000;
        mem[4751] = 12'b011111111000;
        mem[4752] = 12'b011111111000;
        mem[4753] = 12'b011111111000;
        mem[4754] = 12'b011111111000;
        mem[4755] = 12'b011111111000;
        mem[4756] = 12'b011111111001;
        mem[4757] = 12'b011111111001;
        mem[4758] = 12'b011111111001;
        mem[4759] = 12'b011111111001;
        mem[4760] = 12'b011111111001;
        mem[4761] = 12'b011111111001;
        mem[4762] = 12'b011111111001;
        mem[4763] = 12'b011111111001;
        mem[4764] = 12'b011111111001;
        mem[4765] = 12'b011111111001;
        mem[4766] = 12'b011111111001;
        mem[4767] = 12'b011111111001;
        mem[4768] = 12'b011111111001;
        mem[4769] = 12'b011111111001;
        mem[4770] = 12'b011111111001;
        mem[4771] = 12'b011111111001;
        mem[4772] = 12'b011111111001;
        mem[4773] = 12'b011111111001;
        mem[4774] = 12'b011111111001;
        mem[4775] = 12'b011111111001;
        mem[4776] = 12'b011111111001;
        mem[4777] = 12'b011111111010;
        mem[4778] = 12'b011111111010;
        mem[4779] = 12'b011111111010;
        mem[4780] = 12'b011111111010;
        mem[4781] = 12'b011111111010;
        mem[4782] = 12'b011111111010;
        mem[4783] = 12'b011111111010;
        mem[4784] = 12'b011111111010;
        mem[4785] = 12'b011111111010;
        mem[4786] = 12'b011111111010;
        mem[4787] = 12'b011111111010;
        mem[4788] = 12'b011111111010;
        mem[4789] = 12'b011111111010;
        mem[4790] = 12'b011111111010;
        mem[4791] = 12'b011111111010;
        mem[4792] = 12'b011111111010;
        mem[4793] = 12'b011111111010;
        mem[4794] = 12'b011111111010;
        mem[4795] = 12'b011111111010;
        mem[4796] = 12'b011111111010;
        mem[4797] = 12'b011111111010;
        mem[4798] = 12'b011111111010;
        mem[4799] = 12'b011111111010;
        mem[4800] = 12'b011111111010;
        mem[4801] = 12'b011111111011;
        mem[4802] = 12'b011111111011;
        mem[4803] = 12'b011111111011;
        mem[4804] = 12'b011111111011;
        mem[4805] = 12'b011111111011;
        mem[4806] = 12'b011111111011;
        mem[4807] = 12'b011111111011;
        mem[4808] = 12'b011111111011;
        mem[4809] = 12'b011111111011;
        mem[4810] = 12'b011111111011;
        mem[4811] = 12'b011111111011;
        mem[4812] = 12'b011111111011;
        mem[4813] = 12'b011111111011;
        mem[4814] = 12'b011111111011;
        mem[4815] = 12'b011111111011;
        mem[4816] = 12'b011111111011;
        mem[4817] = 12'b011111111011;
        mem[4818] = 12'b011111111011;
        mem[4819] = 12'b011111111011;
        mem[4820] = 12'b011111111011;
        mem[4821] = 12'b011111111011;
        mem[4822] = 12'b011111111011;
        mem[4823] = 12'b011111111011;
        mem[4824] = 12'b011111111011;
        mem[4825] = 12'b011111111011;
        mem[4826] = 12'b011111111011;
        mem[4827] = 12'b011111111011;
        mem[4828] = 12'b011111111100;
        mem[4829] = 12'b011111111100;
        mem[4830] = 12'b011111111100;
        mem[4831] = 12'b011111111100;
        mem[4832] = 12'b011111111100;
        mem[4833] = 12'b011111111100;
        mem[4834] = 12'b011111111100;
        mem[4835] = 12'b011111111100;
        mem[4836] = 12'b011111111100;
        mem[4837] = 12'b011111111100;
        mem[4838] = 12'b011111111100;
        mem[4839] = 12'b011111111100;
        mem[4840] = 12'b011111111100;
        mem[4841] = 12'b011111111100;
        mem[4842] = 12'b011111111100;
        mem[4843] = 12'b011111111100;
        mem[4844] = 12'b011111111100;
        mem[4845] = 12'b011111111100;
        mem[4846] = 12'b011111111100;
        mem[4847] = 12'b011111111100;
        mem[4848] = 12'b011111111100;
        mem[4849] = 12'b011111111100;
        mem[4850] = 12'b011111111100;
        mem[4851] = 12'b011111111100;
        mem[4852] = 12'b011111111100;
        mem[4853] = 12'b011111111100;
        mem[4854] = 12'b011111111100;
        mem[4855] = 12'b011111111100;
        mem[4856] = 12'b011111111100;
        mem[4857] = 12'b011111111100;
        mem[4858] = 12'b011111111100;
        mem[4859] = 12'b011111111101;
        mem[4860] = 12'b011111111101;
        mem[4861] = 12'b011111111101;
        mem[4862] = 12'b011111111101;
        mem[4863] = 12'b011111111101;
        mem[4864] = 12'b011111111101;
        mem[4865] = 12'b011111111101;
        mem[4866] = 12'b011111111101;
        mem[4867] = 12'b011111111101;
        mem[4868] = 12'b011111111101;
        mem[4869] = 12'b011111111101;
        mem[4870] = 12'b011111111101;
        mem[4871] = 12'b011111111101;
        mem[4872] = 12'b011111111101;
        mem[4873] = 12'b011111111101;
        mem[4874] = 12'b011111111101;
        mem[4875] = 12'b011111111101;
        mem[4876] = 12'b011111111101;
        mem[4877] = 12'b011111111101;
        mem[4878] = 12'b011111111101;
        mem[4879] = 12'b011111111101;
        mem[4880] = 12'b011111111101;
        mem[4881] = 12'b011111111101;
        mem[4882] = 12'b011111111101;
        mem[4883] = 12'b011111111101;
        mem[4884] = 12'b011111111101;
        mem[4885] = 12'b011111111101;
        mem[4886] = 12'b011111111101;
        mem[4887] = 12'b011111111101;
        mem[4888] = 12'b011111111101;
        mem[4889] = 12'b011111111101;
        mem[4890] = 12'b011111111101;
        mem[4891] = 12'b011111111101;
        mem[4892] = 12'b011111111101;
        mem[4893] = 12'b011111111101;
        mem[4894] = 12'b011111111101;
        mem[4895] = 12'b011111111101;
        mem[4896] = 12'b011111111101;
        mem[4897] = 12'b011111111101;
        mem[4898] = 12'b011111111101;
        mem[4899] = 12'b011111111101;
        mem[4900] = 12'b011111111101;
        mem[4901] = 12'b011111111110;
        mem[4902] = 12'b011111111110;
        mem[4903] = 12'b011111111110;
        mem[4904] = 12'b011111111110;
        mem[4905] = 12'b011111111110;
        mem[4906] = 12'b011111111110;
        mem[4907] = 12'b011111111110;
        mem[4908] = 12'b011111111110;
        mem[4909] = 12'b011111111110;
        mem[4910] = 12'b011111111110;
        mem[4911] = 12'b011111111110;
        mem[4912] = 12'b011111111110;
        mem[4913] = 12'b011111111110;
        mem[4914] = 12'b011111111110;
        mem[4915] = 12'b011111111110;
        mem[4916] = 12'b011111111110;
        mem[4917] = 12'b011111111110;
        mem[4918] = 12'b011111111110;
        mem[4919] = 12'b011111111110;
        mem[4920] = 12'b011111111110;
        mem[4921] = 12'b011111111110;
        mem[4922] = 12'b011111111110;
        mem[4923] = 12'b011111111110;
        mem[4924] = 12'b011111111110;
        mem[4925] = 12'b011111111110;
        mem[4926] = 12'b011111111110;
        mem[4927] = 12'b011111111110;
        mem[4928] = 12'b011111111110;
        mem[4929] = 12'b011111111110;
        mem[4930] = 12'b011111111110;
        mem[4931] = 12'b011111111110;
        mem[4932] = 12'b011111111110;
        mem[4933] = 12'b011111111110;
        mem[4934] = 12'b011111111110;
        mem[4935] = 12'b011111111110;
        mem[4936] = 12'b011111111110;
        mem[4937] = 12'b011111111110;
        mem[4938] = 12'b011111111110;
        mem[4939] = 12'b011111111110;
        mem[4940] = 12'b011111111110;
        mem[4941] = 12'b011111111110;
        mem[4942] = 12'b011111111110;
        mem[4943] = 12'b011111111110;
        mem[4944] = 12'b011111111110;
        mem[4945] = 12'b011111111110;
        mem[4946] = 12'b011111111110;
        mem[4947] = 12'b011111111110;
        mem[4948] = 12'b011111111110;
        mem[4949] = 12'b011111111110;
        mem[4950] = 12'b011111111110;
        mem[4951] = 12'b011111111110;
        mem[4952] = 12'b011111111110;
        mem[4953] = 12'b011111111110;
        mem[4954] = 12'b011111111110;
        mem[4955] = 12'b011111111110;
        mem[4956] = 12'b011111111110;
        mem[4957] = 12'b011111111110;
        mem[4958] = 12'b011111111110;
        mem[4959] = 12'b011111111110;
        mem[4960] = 12'b011111111110;
        mem[4961] = 12'b011111111110;
        mem[4962] = 12'b011111111110;
        mem[4963] = 12'b011111111110;
        mem[4964] = 12'b011111111110;
        mem[4965] = 12'b011111111110;
        mem[4966] = 12'b011111111110;
        mem[4967] = 12'b011111111110;
        mem[4968] = 12'b011111111110;
        mem[4969] = 12'b011111111110;
        mem[4970] = 12'b011111111110;
        mem[4971] = 12'b011111111110;
        mem[4972] = 12'b011111111110;
        mem[4973] = 12'b011111111110;
        mem[4974] = 12'b011111111110;
        mem[4975] = 12'b011111111110;
        mem[4976] = 12'b011111111110;
        mem[4977] = 12'b011111111110;
        mem[4978] = 12'b011111111110;
        mem[4979] = 12'b011111111110;
        mem[4980] = 12'b011111111110;
        mem[4981] = 12'b011111111110;
        mem[4982] = 12'b011111111110;
        mem[4983] = 12'b011111111110;
        mem[4984] = 12'b011111111110;
        mem[4985] = 12'b011111111110;
        mem[4986] = 12'b011111111110;
        mem[4987] = 12'b011111111110;
        mem[4988] = 12'b011111111110;
        mem[4989] = 12'b011111111110;
        mem[4990] = 12'b011111111110;
        mem[4991] = 12'b011111111110;
        mem[4992] = 12'b011111111110;
        mem[4993] = 12'b011111111110;
        mem[4994] = 12'b011111111110;
        mem[4995] = 12'b011111111110;
        mem[4996] = 12'b011111111110;
        mem[4997] = 12'b011111111110;
        mem[4998] = 12'b011111111110;
        mem[4999] = 12'b011111111110;
        mem[5000] = 12'b011111111110;
        mem[5001] = 12'b011111111110;
        mem[5002] = 12'b011111111110;
        mem[5003] = 12'b011111111110;
        mem[5004] = 12'b011111111110;
        mem[5005] = 12'b011111111110;
        mem[5006] = 12'b011111111110;
        mem[5007] = 12'b011111111110;
        mem[5008] = 12'b011111111110;
        mem[5009] = 12'b011111111110;
        mem[5010] = 12'b011111111110;
        mem[5011] = 12'b011111111110;
        mem[5012] = 12'b011111111110;
        mem[5013] = 12'b011111111110;
        mem[5014] = 12'b011111111110;
        mem[5015] = 12'b011111111110;
        mem[5016] = 12'b011111111110;
        mem[5017] = 12'b011111111110;
        mem[5018] = 12'b011111111110;
        mem[5019] = 12'b011111111110;
        mem[5020] = 12'b011111111110;
        mem[5021] = 12'b011111111110;
        mem[5022] = 12'b011111111110;
        mem[5023] = 12'b011111111110;
        mem[5024] = 12'b011111111110;
        mem[5025] = 12'b011111111110;
        mem[5026] = 12'b011111111110;
        mem[5027] = 12'b011111111110;
        mem[5028] = 12'b011111111110;
        mem[5029] = 12'b011111111110;
        mem[5030] = 12'b011111111110;
        mem[5031] = 12'b011111111110;
        mem[5032] = 12'b011111111110;
        mem[5033] = 12'b011111111110;
        mem[5034] = 12'b011111111110;
        mem[5035] = 12'b011111111110;
        mem[5036] = 12'b011111111110;
        mem[5037] = 12'b011111111110;
        mem[5038] = 12'b011111111110;
        mem[5039] = 12'b011111111110;
        mem[5040] = 12'b011111111110;
        mem[5041] = 12'b011111111110;
        mem[5042] = 12'b011111111110;
        mem[5043] = 12'b011111111110;
        mem[5044] = 12'b011111111110;
        mem[5045] = 12'b011111111110;
        mem[5046] = 12'b011111111110;
        mem[5047] = 12'b011111111110;
        mem[5048] = 12'b011111111110;
        mem[5049] = 12'b011111111110;
        mem[5050] = 12'b011111111110;
        mem[5051] = 12'b011111111110;
        mem[5052] = 12'b011111111110;
        mem[5053] = 12'b011111111110;
        mem[5054] = 12'b011111111110;
        mem[5055] = 12'b011111111110;
        mem[5056] = 12'b011111111110;
        mem[5057] = 12'b011111111110;
        mem[5058] = 12'b011111111110;
        mem[5059] = 12'b011111111110;
        mem[5060] = 12'b011111111110;
        mem[5061] = 12'b011111111110;
        mem[5062] = 12'b011111111110;
        mem[5063] = 12'b011111111110;
        mem[5064] = 12'b011111111110;
        mem[5065] = 12'b011111111110;
        mem[5066] = 12'b011111111110;
        mem[5067] = 12'b011111111110;
        mem[5068] = 12'b011111111110;
        mem[5069] = 12'b011111111110;
        mem[5070] = 12'b011111111110;
        mem[5071] = 12'b011111111110;
        mem[5072] = 12'b011111111110;
        mem[5073] = 12'b011111111110;
        mem[5074] = 12'b011111111110;
        mem[5075] = 12'b011111111110;
        mem[5076] = 12'b011111111110;
        mem[5077] = 12'b011111111110;
        mem[5078] = 12'b011111111110;
        mem[5079] = 12'b011111111110;
        mem[5080] = 12'b011111111110;
        mem[5081] = 12'b011111111110;
        mem[5082] = 12'b011111111110;
        mem[5083] = 12'b011111111110;
        mem[5084] = 12'b011111111110;
        mem[5085] = 12'b011111111110;
        mem[5086] = 12'b011111111110;
        mem[5087] = 12'b011111111110;
        mem[5088] = 12'b011111111110;
        mem[5089] = 12'b011111111110;
        mem[5090] = 12'b011111111110;
        mem[5091] = 12'b011111111110;
        mem[5092] = 12'b011111111110;
        mem[5093] = 12'b011111111110;
        mem[5094] = 12'b011111111110;
        mem[5095] = 12'b011111111110;
        mem[5096] = 12'b011111111110;
        mem[5097] = 12'b011111111110;
        mem[5098] = 12'b011111111110;
        mem[5099] = 12'b011111111101;
        mem[5100] = 12'b011111111101;
        mem[5101] = 12'b011111111101;
        mem[5102] = 12'b011111111101;
        mem[5103] = 12'b011111111101;
        mem[5104] = 12'b011111111101;
        mem[5105] = 12'b011111111101;
        mem[5106] = 12'b011111111101;
        mem[5107] = 12'b011111111101;
        mem[5108] = 12'b011111111101;
        mem[5109] = 12'b011111111101;
        mem[5110] = 12'b011111111101;
        mem[5111] = 12'b011111111101;
        mem[5112] = 12'b011111111101;
        mem[5113] = 12'b011111111101;
        mem[5114] = 12'b011111111101;
        mem[5115] = 12'b011111111101;
        mem[5116] = 12'b011111111101;
        mem[5117] = 12'b011111111101;
        mem[5118] = 12'b011111111101;
        mem[5119] = 12'b011111111101;
        mem[5120] = 12'b011111111101;
        mem[5121] = 12'b011111111101;
        mem[5122] = 12'b011111111101;
        mem[5123] = 12'b011111111101;
        mem[5124] = 12'b011111111101;
        mem[5125] = 12'b011111111101;
        mem[5126] = 12'b011111111101;
        mem[5127] = 12'b011111111101;
        mem[5128] = 12'b011111111101;
        mem[5129] = 12'b011111111101;
        mem[5130] = 12'b011111111101;
        mem[5131] = 12'b011111111101;
        mem[5132] = 12'b011111111101;
        mem[5133] = 12'b011111111101;
        mem[5134] = 12'b011111111101;
        mem[5135] = 12'b011111111101;
        mem[5136] = 12'b011111111101;
        mem[5137] = 12'b011111111101;
        mem[5138] = 12'b011111111101;
        mem[5139] = 12'b011111111101;
        mem[5140] = 12'b011111111101;
        mem[5141] = 12'b011111111100;
        mem[5142] = 12'b011111111100;
        mem[5143] = 12'b011111111100;
        mem[5144] = 12'b011111111100;
        mem[5145] = 12'b011111111100;
        mem[5146] = 12'b011111111100;
        mem[5147] = 12'b011111111100;
        mem[5148] = 12'b011111111100;
        mem[5149] = 12'b011111111100;
        mem[5150] = 12'b011111111100;
        mem[5151] = 12'b011111111100;
        mem[5152] = 12'b011111111100;
        mem[5153] = 12'b011111111100;
        mem[5154] = 12'b011111111100;
        mem[5155] = 12'b011111111100;
        mem[5156] = 12'b011111111100;
        mem[5157] = 12'b011111111100;
        mem[5158] = 12'b011111111100;
        mem[5159] = 12'b011111111100;
        mem[5160] = 12'b011111111100;
        mem[5161] = 12'b011111111100;
        mem[5162] = 12'b011111111100;
        mem[5163] = 12'b011111111100;
        mem[5164] = 12'b011111111100;
        mem[5165] = 12'b011111111100;
        mem[5166] = 12'b011111111100;
        mem[5167] = 12'b011111111100;
        mem[5168] = 12'b011111111100;
        mem[5169] = 12'b011111111100;
        mem[5170] = 12'b011111111100;
        mem[5171] = 12'b011111111100;
        mem[5172] = 12'b011111111011;
        mem[5173] = 12'b011111111011;
        mem[5174] = 12'b011111111011;
        mem[5175] = 12'b011111111011;
        mem[5176] = 12'b011111111011;
        mem[5177] = 12'b011111111011;
        mem[5178] = 12'b011111111011;
        mem[5179] = 12'b011111111011;
        mem[5180] = 12'b011111111011;
        mem[5181] = 12'b011111111011;
        mem[5182] = 12'b011111111011;
        mem[5183] = 12'b011111111011;
        mem[5184] = 12'b011111111011;
        mem[5185] = 12'b011111111011;
        mem[5186] = 12'b011111111011;
        mem[5187] = 12'b011111111011;
        mem[5188] = 12'b011111111011;
        mem[5189] = 12'b011111111011;
        mem[5190] = 12'b011111111011;
        mem[5191] = 12'b011111111011;
        mem[5192] = 12'b011111111011;
        mem[5193] = 12'b011111111011;
        mem[5194] = 12'b011111111011;
        mem[5195] = 12'b011111111011;
        mem[5196] = 12'b011111111011;
        mem[5197] = 12'b011111111011;
        mem[5198] = 12'b011111111011;
        mem[5199] = 12'b011111111010;
        mem[5200] = 12'b011111111010;
        mem[5201] = 12'b011111111010;
        mem[5202] = 12'b011111111010;
        mem[5203] = 12'b011111111010;
        mem[5204] = 12'b011111111010;
        mem[5205] = 12'b011111111010;
        mem[5206] = 12'b011111111010;
        mem[5207] = 12'b011111111010;
        mem[5208] = 12'b011111111010;
        mem[5209] = 12'b011111111010;
        mem[5210] = 12'b011111111010;
        mem[5211] = 12'b011111111010;
        mem[5212] = 12'b011111111010;
        mem[5213] = 12'b011111111010;
        mem[5214] = 12'b011111111010;
        mem[5215] = 12'b011111111010;
        mem[5216] = 12'b011111111010;
        mem[5217] = 12'b011111111010;
        mem[5218] = 12'b011111111010;
        mem[5219] = 12'b011111111010;
        mem[5220] = 12'b011111111010;
        mem[5221] = 12'b011111111010;
        mem[5222] = 12'b011111111010;
        mem[5223] = 12'b011111111001;
        mem[5224] = 12'b011111111001;
        mem[5225] = 12'b011111111001;
        mem[5226] = 12'b011111111001;
        mem[5227] = 12'b011111111001;
        mem[5228] = 12'b011111111001;
        mem[5229] = 12'b011111111001;
        mem[5230] = 12'b011111111001;
        mem[5231] = 12'b011111111001;
        mem[5232] = 12'b011111111001;
        mem[5233] = 12'b011111111001;
        mem[5234] = 12'b011111111001;
        mem[5235] = 12'b011111111001;
        mem[5236] = 12'b011111111001;
        mem[5237] = 12'b011111111001;
        mem[5238] = 12'b011111111001;
        mem[5239] = 12'b011111111001;
        mem[5240] = 12'b011111111001;
        mem[5241] = 12'b011111111001;
        mem[5242] = 12'b011111111001;
        mem[5243] = 12'b011111111001;
        mem[5244] = 12'b011111111000;
        mem[5245] = 12'b011111111000;
        mem[5246] = 12'b011111111000;
        mem[5247] = 12'b011111111000;
        mem[5248] = 12'b011111111000;
        mem[5249] = 12'b011111111000;
        mem[5250] = 12'b011111111000;
        mem[5251] = 12'b011111111000;
        mem[5252] = 12'b011111111000;
        mem[5253] = 12'b011111111000;
        mem[5254] = 12'b011111111000;
        mem[5255] = 12'b011111111000;
        mem[5256] = 12'b011111111000;
        mem[5257] = 12'b011111111000;
        mem[5258] = 12'b011111111000;
        mem[5259] = 12'b011111111000;
        mem[5260] = 12'b011111111000;
        mem[5261] = 12'b011111111000;
        mem[5262] = 12'b011111111000;
        mem[5263] = 12'b011111110111;
        mem[5264] = 12'b011111110111;
        mem[5265] = 12'b011111110111;
        mem[5266] = 12'b011111110111;
        mem[5267] = 12'b011111110111;
        mem[5268] = 12'b011111110111;
        mem[5269] = 12'b011111110111;
        mem[5270] = 12'b011111110111;
        mem[5271] = 12'b011111110111;
        mem[5272] = 12'b011111110111;
        mem[5273] = 12'b011111110111;
        mem[5274] = 12'b011111110111;
        mem[5275] = 12'b011111110111;
        mem[5276] = 12'b011111110111;
        mem[5277] = 12'b011111110111;
        mem[5278] = 12'b011111110111;
        mem[5279] = 12'b011111110111;
        mem[5280] = 12'b011111110111;
        mem[5281] = 12'b011111110110;
        mem[5282] = 12'b011111110110;
        mem[5283] = 12'b011111110110;
        mem[5284] = 12'b011111110110;
        mem[5285] = 12'b011111110110;
        mem[5286] = 12'b011111110110;
        mem[5287] = 12'b011111110110;
        mem[5288] = 12'b011111110110;
        mem[5289] = 12'b011111110110;
        mem[5290] = 12'b011111110110;
        mem[5291] = 12'b011111110110;
        mem[5292] = 12'b011111110110;
        mem[5293] = 12'b011111110110;
        mem[5294] = 12'b011111110110;
        mem[5295] = 12'b011111110110;
        mem[5296] = 12'b011111110110;
        mem[5297] = 12'b011111110110;
        mem[5298] = 12'b011111110110;
        mem[5299] = 12'b011111110101;
        mem[5300] = 12'b011111110101;
        mem[5301] = 12'b011111110101;
        mem[5302] = 12'b011111110101;
        mem[5303] = 12'b011111110101;
        mem[5304] = 12'b011111110101;
        mem[5305] = 12'b011111110101;
        mem[5306] = 12'b011111110101;
        mem[5307] = 12'b011111110101;
        mem[5308] = 12'b011111110101;
        mem[5309] = 12'b011111110101;
        mem[5310] = 12'b011111110101;
        mem[5311] = 12'b011111110101;
        mem[5312] = 12'b011111110101;
        mem[5313] = 12'b011111110101;
        mem[5314] = 12'b011111110101;
        mem[5315] = 12'b011111110100;
        mem[5316] = 12'b011111110100;
        mem[5317] = 12'b011111110100;
        mem[5318] = 12'b011111110100;
        mem[5319] = 12'b011111110100;
        mem[5320] = 12'b011111110100;
        mem[5321] = 12'b011111110100;
        mem[5322] = 12'b011111110100;
        mem[5323] = 12'b011111110100;
        mem[5324] = 12'b011111110100;
        mem[5325] = 12'b011111110100;
        mem[5326] = 12'b011111110100;
        mem[5327] = 12'b011111110100;
        mem[5328] = 12'b011111110100;
        mem[5329] = 12'b011111110100;
        mem[5330] = 12'b011111110011;
        mem[5331] = 12'b011111110011;
        mem[5332] = 12'b011111110011;
        mem[5333] = 12'b011111110011;
        mem[5334] = 12'b011111110011;
        mem[5335] = 12'b011111110011;
        mem[5336] = 12'b011111110011;
        mem[5337] = 12'b011111110011;
        mem[5338] = 12'b011111110011;
        mem[5339] = 12'b011111110011;
        mem[5340] = 12'b011111110011;
        mem[5341] = 12'b011111110011;
        mem[5342] = 12'b011111110011;
        mem[5343] = 12'b011111110011;
        mem[5344] = 12'b011111110011;
        mem[5345] = 12'b011111110010;
        mem[5346] = 12'b011111110010;
        mem[5347] = 12'b011111110010;
        mem[5348] = 12'b011111110010;
        mem[5349] = 12'b011111110010;
        mem[5350] = 12'b011111110010;
        mem[5351] = 12'b011111110010;
        mem[5352] = 12'b011111110010;
        mem[5353] = 12'b011111110010;
        mem[5354] = 12'b011111110010;
        mem[5355] = 12'b011111110010;
        mem[5356] = 12'b011111110010;
        mem[5357] = 12'b011111110010;
        mem[5358] = 12'b011111110010;
        mem[5359] = 12'b011111110001;
        mem[5360] = 12'b011111110001;
        mem[5361] = 12'b011111110001;
        mem[5362] = 12'b011111110001;
        mem[5363] = 12'b011111110001;
        mem[5364] = 12'b011111110001;
        mem[5365] = 12'b011111110001;
        mem[5366] = 12'b011111110001;
        mem[5367] = 12'b011111110001;
        mem[5368] = 12'b011111110001;
        mem[5369] = 12'b011111110001;
        mem[5370] = 12'b011111110001;
        mem[5371] = 12'b011111110001;
        mem[5372] = 12'b011111110000;
        mem[5373] = 12'b011111110000;
        mem[5374] = 12'b011111110000;
        mem[5375] = 12'b011111110000;
        mem[5376] = 12'b011111110000;
        mem[5377] = 12'b011111110000;
        mem[5378] = 12'b011111110000;
        mem[5379] = 12'b011111110000;
        mem[5380] = 12'b011111110000;
        mem[5381] = 12'b011111110000;
        mem[5382] = 12'b011111110000;
        mem[5383] = 12'b011111110000;
        mem[5384] = 12'b011111110000;
        mem[5385] = 12'b011111110000;
        mem[5386] = 12'b011111101111;
        mem[5387] = 12'b011111101111;
        mem[5388] = 12'b011111101111;
        mem[5389] = 12'b011111101111;
        mem[5390] = 12'b011111101111;
        mem[5391] = 12'b011111101111;
        mem[5392] = 12'b011111101111;
        mem[5393] = 12'b011111101111;
        mem[5394] = 12'b011111101111;
        mem[5395] = 12'b011111101111;
        mem[5396] = 12'b011111101111;
        mem[5397] = 12'b011111101111;
        mem[5398] = 12'b011111101110;
        mem[5399] = 12'b011111101110;
        mem[5400] = 12'b011111101110;
        mem[5401] = 12'b011111101110;
        mem[5402] = 12'b011111101110;
        mem[5403] = 12'b011111101110;
        mem[5404] = 12'b011111101110;
        mem[5405] = 12'b011111101110;
        mem[5406] = 12'b011111101110;
        mem[5407] = 12'b011111101110;
        mem[5408] = 12'b011111101110;
        mem[5409] = 12'b011111101110;
        mem[5410] = 12'b011111101101;
        mem[5411] = 12'b011111101101;
        mem[5412] = 12'b011111101101;
        mem[5413] = 12'b011111101101;
        mem[5414] = 12'b011111101101;
        mem[5415] = 12'b011111101101;
        mem[5416] = 12'b011111101101;
        mem[5417] = 12'b011111101101;
        mem[5418] = 12'b011111101101;
        mem[5419] = 12'b011111101101;
        mem[5420] = 12'b011111101101;
        mem[5421] = 12'b011111101101;
        mem[5422] = 12'b011111101100;
        mem[5423] = 12'b011111101100;
        mem[5424] = 12'b011111101100;
        mem[5425] = 12'b011111101100;
        mem[5426] = 12'b011111101100;
        mem[5427] = 12'b011111101100;
        mem[5428] = 12'b011111101100;
        mem[5429] = 12'b011111101100;
        mem[5430] = 12'b011111101100;
        mem[5431] = 12'b011111101100;
        mem[5432] = 12'b011111101100;
        mem[5433] = 12'b011111101100;
        mem[5434] = 12'b011111101011;
        mem[5435] = 12'b011111101011;
        mem[5436] = 12'b011111101011;
        mem[5437] = 12'b011111101011;
        mem[5438] = 12'b011111101011;
        mem[5439] = 12'b011111101011;
        mem[5440] = 12'b011111101011;
        mem[5441] = 12'b011111101011;
        mem[5442] = 12'b011111101011;
        mem[5443] = 12'b011111101011;
        mem[5444] = 12'b011111101011;
        mem[5445] = 12'b011111101010;
        mem[5446] = 12'b011111101010;
        mem[5447] = 12'b011111101010;
        mem[5448] = 12'b011111101010;
        mem[5449] = 12'b011111101010;
        mem[5450] = 12'b011111101010;
        mem[5451] = 12'b011111101010;
        mem[5452] = 12'b011111101010;
        mem[5453] = 12'b011111101010;
        mem[5454] = 12'b011111101010;
        mem[5455] = 12'b011111101010;
        mem[5456] = 12'b011111101001;
        mem[5457] = 12'b011111101001;
        mem[5458] = 12'b011111101001;
        mem[5459] = 12'b011111101001;
        mem[5460] = 12'b011111101001;
        mem[5461] = 12'b011111101001;
        mem[5462] = 12'b011111101001;
        mem[5463] = 12'b011111101001;
        mem[5464] = 12'b011111101001;
        mem[5465] = 12'b011111101001;
        mem[5466] = 12'b011111101001;
        mem[5467] = 12'b011111101000;
        mem[5468] = 12'b011111101000;
        mem[5469] = 12'b011111101000;
        mem[5470] = 12'b011111101000;
        mem[5471] = 12'b011111101000;
        mem[5472] = 12'b011111101000;
        mem[5473] = 12'b011111101000;
        mem[5474] = 12'b011111101000;
        mem[5475] = 12'b011111101000;
        mem[5476] = 12'b011111101000;
        mem[5477] = 12'b011111101000;
        mem[5478] = 12'b011111100111;
        mem[5479] = 12'b011111100111;
        mem[5480] = 12'b011111100111;
        mem[5481] = 12'b011111100111;
        mem[5482] = 12'b011111100111;
        mem[5483] = 12'b011111100111;
        mem[5484] = 12'b011111100111;
        mem[5485] = 12'b011111100111;
        mem[5486] = 12'b011111100111;
        mem[5487] = 12'b011111100111;
        mem[5488] = 12'b011111100110;
        mem[5489] = 12'b011111100110;
        mem[5490] = 12'b011111100110;
        mem[5491] = 12'b011111100110;
        mem[5492] = 12'b011111100110;
        mem[5493] = 12'b011111100110;
        mem[5494] = 12'b011111100110;
        mem[5495] = 12'b011111100110;
        mem[5496] = 12'b011111100110;
        mem[5497] = 12'b011111100110;
        mem[5498] = 12'b011111100101;
        mem[5499] = 12'b011111100101;
        mem[5500] = 12'b011111100101;
        mem[5501] = 12'b011111100101;
        mem[5502] = 12'b011111100101;
        mem[5503] = 12'b011111100101;
        mem[5504] = 12'b011111100101;
        mem[5505] = 12'b011111100101;
        mem[5506] = 12'b011111100101;
        mem[5507] = 12'b011111100101;
        mem[5508] = 12'b011111100100;
        mem[5509] = 12'b011111100100;
        mem[5510] = 12'b011111100100;
        mem[5511] = 12'b011111100100;
        mem[5512] = 12'b011111100100;
        mem[5513] = 12'b011111100100;
        mem[5514] = 12'b011111100100;
        mem[5515] = 12'b011111100100;
        mem[5516] = 12'b011111100100;
        mem[5517] = 12'b011111100100;
        mem[5518] = 12'b011111100011;
        mem[5519] = 12'b011111100011;
        mem[5520] = 12'b011111100011;
        mem[5521] = 12'b011111100011;
        mem[5522] = 12'b011111100011;
        mem[5523] = 12'b011111100011;
        mem[5524] = 12'b011111100011;
        mem[5525] = 12'b011111100011;
        mem[5526] = 12'b011111100011;
        mem[5527] = 12'b011111100010;
        mem[5528] = 12'b011111100010;
        mem[5529] = 12'b011111100010;
        mem[5530] = 12'b011111100010;
        mem[5531] = 12'b011111100010;
        mem[5532] = 12'b011111100010;
        mem[5533] = 12'b011111100010;
        mem[5534] = 12'b011111100010;
        mem[5535] = 12'b011111100010;
        mem[5536] = 12'b011111100001;
        mem[5537] = 12'b011111100001;
        mem[5538] = 12'b011111100001;
        mem[5539] = 12'b011111100001;
        mem[5540] = 12'b011111100001;
        mem[5541] = 12'b011111100001;
        mem[5542] = 12'b011111100001;
        mem[5543] = 12'b011111100001;
        mem[5544] = 12'b011111100001;
        mem[5545] = 12'b011111100001;
        mem[5546] = 12'b011111100000;
        mem[5547] = 12'b011111100000;
        mem[5548] = 12'b011111100000;
        mem[5549] = 12'b011111100000;
        mem[5550] = 12'b011111100000;
        mem[5551] = 12'b011111100000;
        mem[5552] = 12'b011111100000;
        mem[5553] = 12'b011111100000;
        mem[5554] = 12'b011111100000;
        mem[5555] = 12'b011111011111;
        mem[5556] = 12'b011111011111;
        mem[5557] = 12'b011111011111;
        mem[5558] = 12'b011111011111;
        mem[5559] = 12'b011111011111;
        mem[5560] = 12'b011111011111;
        mem[5561] = 12'b011111011111;
        mem[5562] = 12'b011111011111;
        mem[5563] = 12'b011111011111;
        mem[5564] = 12'b011111011110;
        mem[5565] = 12'b011111011110;
        mem[5566] = 12'b011111011110;
        mem[5567] = 12'b011111011110;
        mem[5568] = 12'b011111011110;
        mem[5569] = 12'b011111011110;
        mem[5570] = 12'b011111011110;
        mem[5571] = 12'b011111011110;
        mem[5572] = 12'b011111011101;
        mem[5573] = 12'b011111011101;
        mem[5574] = 12'b011111011101;
        mem[5575] = 12'b011111011101;
        mem[5576] = 12'b011111011101;
        mem[5577] = 12'b011111011101;
        mem[5578] = 12'b011111011101;
        mem[5579] = 12'b011111011101;
        mem[5580] = 12'b011111011101;
        mem[5581] = 12'b011111011100;
        mem[5582] = 12'b011111011100;
        mem[5583] = 12'b011111011100;
        mem[5584] = 12'b011111011100;
        mem[5585] = 12'b011111011100;
        mem[5586] = 12'b011111011100;
        mem[5587] = 12'b011111011100;
        mem[5588] = 12'b011111011100;
        mem[5589] = 12'b011111011011;
        mem[5590] = 12'b011111011011;
        mem[5591] = 12'b011111011011;
        mem[5592] = 12'b011111011011;
        mem[5593] = 12'b011111011011;
        mem[5594] = 12'b011111011011;
        mem[5595] = 12'b011111011011;
        mem[5596] = 12'b011111011011;
        mem[5597] = 12'b011111011011;
        mem[5598] = 12'b011111011010;
        mem[5599] = 12'b011111011010;
        mem[5600] = 12'b011111011010;
        mem[5601] = 12'b011111011010;
        mem[5602] = 12'b011111011010;
        mem[5603] = 12'b011111011010;
        mem[5604] = 12'b011111011010;
        mem[5605] = 12'b011111011010;
        mem[5606] = 12'b011111011001;
        mem[5607] = 12'b011111011001;
        mem[5608] = 12'b011111011001;
        mem[5609] = 12'b011111011001;
        mem[5610] = 12'b011111011001;
        mem[5611] = 12'b011111011001;
        mem[5612] = 12'b011111011001;
        mem[5613] = 12'b011111011001;
        mem[5614] = 12'b011111011000;
        mem[5615] = 12'b011111011000;
        mem[5616] = 12'b011111011000;
        mem[5617] = 12'b011111011000;
        mem[5618] = 12'b011111011000;
        mem[5619] = 12'b011111011000;
        mem[5620] = 12'b011111011000;
        mem[5621] = 12'b011111011000;
        mem[5622] = 12'b011111010111;
        mem[5623] = 12'b011111010111;
        mem[5624] = 12'b011111010111;
        mem[5625] = 12'b011111010111;
        mem[5626] = 12'b011111010111;
        mem[5627] = 12'b011111010111;
        mem[5628] = 12'b011111010111;
        mem[5629] = 12'b011111010111;
        mem[5630] = 12'b011111010110;
        mem[5631] = 12'b011111010110;
        mem[5632] = 12'b011111010110;
        mem[5633] = 12'b011111010110;
        mem[5634] = 12'b011111010110;
        mem[5635] = 12'b011111010110;
        mem[5636] = 12'b011111010110;
        mem[5637] = 12'b011111010110;
        mem[5638] = 12'b011111010101;
        mem[5639] = 12'b011111010101;
        mem[5640] = 12'b011111010101;
        mem[5641] = 12'b011111010101;
        mem[5642] = 12'b011111010101;
        mem[5643] = 12'b011111010101;
        mem[5644] = 12'b011111010101;
        mem[5645] = 12'b011111010101;
        mem[5646] = 12'b011111010100;
        mem[5647] = 12'b011111010100;
        mem[5648] = 12'b011111010100;
        mem[5649] = 12'b011111010100;
        mem[5650] = 12'b011111010100;
        mem[5651] = 12'b011111010100;
        mem[5652] = 12'b011111010100;
        mem[5653] = 12'b011111010100;
        mem[5654] = 12'b011111010011;
        mem[5655] = 12'b011111010011;
        mem[5656] = 12'b011111010011;
        mem[5657] = 12'b011111010011;
        mem[5658] = 12'b011111010011;
        mem[5659] = 12'b011111010011;
        mem[5660] = 12'b011111010011;
        mem[5661] = 12'b011111010010;
        mem[5662] = 12'b011111010010;
        mem[5663] = 12'b011111010010;
        mem[5664] = 12'b011111010010;
        mem[5665] = 12'b011111010010;
        mem[5666] = 12'b011111010010;
        mem[5667] = 12'b011111010010;
        mem[5668] = 12'b011111010010;
        mem[5669] = 12'b011111010001;
        mem[5670] = 12'b011111010001;
        mem[5671] = 12'b011111010001;
        mem[5672] = 12'b011111010001;
        mem[5673] = 12'b011111010001;
        mem[5674] = 12'b011111010001;
        mem[5675] = 12'b011111010001;
        mem[5676] = 12'b011111010000;
        mem[5677] = 12'b011111010000;
        mem[5678] = 12'b011111010000;
        mem[5679] = 12'b011111010000;
        mem[5680] = 12'b011111010000;
        mem[5681] = 12'b011111010000;
        mem[5682] = 12'b011111010000;
        mem[5683] = 12'b011111001111;
        mem[5684] = 12'b011111001111;
        mem[5685] = 12'b011111001111;
        mem[5686] = 12'b011111001111;
        mem[5687] = 12'b011111001111;
        mem[5688] = 12'b011111001111;
        mem[5689] = 12'b011111001111;
        mem[5690] = 12'b011111001111;
        mem[5691] = 12'b011111001110;
        mem[5692] = 12'b011111001110;
        mem[5693] = 12'b011111001110;
        mem[5694] = 12'b011111001110;
        mem[5695] = 12'b011111001110;
        mem[5696] = 12'b011111001110;
        mem[5697] = 12'b011111001110;
        mem[5698] = 12'b011111001101;
        mem[5699] = 12'b011111001101;
        mem[5700] = 12'b011111001101;
        mem[5701] = 12'b011111001101;
        mem[5702] = 12'b011111001101;
        mem[5703] = 12'b011111001101;
        mem[5704] = 12'b011111001101;
        mem[5705] = 12'b011111001100;
        mem[5706] = 12'b011111001100;
        mem[5707] = 12'b011111001100;
        mem[5708] = 12'b011111001100;
        mem[5709] = 12'b011111001100;
        mem[5710] = 12'b011111001100;
        mem[5711] = 12'b011111001100;
        mem[5712] = 12'b011111001011;
        mem[5713] = 12'b011111001011;
        mem[5714] = 12'b011111001011;
        mem[5715] = 12'b011111001011;
        mem[5716] = 12'b011111001011;
        mem[5717] = 12'b011111001011;
        mem[5718] = 12'b011111001011;
        mem[5719] = 12'b011111001010;
        mem[5720] = 12'b011111001010;
        mem[5721] = 12'b011111001010;
        mem[5722] = 12'b011111001010;
        mem[5723] = 12'b011111001010;
        mem[5724] = 12'b011111001010;
        mem[5725] = 12'b011111001010;
        mem[5726] = 12'b011111001001;
        mem[5727] = 12'b011111001001;
        mem[5728] = 12'b011111001001;
        mem[5729] = 12'b011111001001;
        mem[5730] = 12'b011111001001;
        mem[5731] = 12'b011111001001;
        mem[5732] = 12'b011111001001;
        mem[5733] = 12'b011111001000;
        mem[5734] = 12'b011111001000;
        mem[5735] = 12'b011111001000;
        mem[5736] = 12'b011111001000;
        mem[5737] = 12'b011111001000;
        mem[5738] = 12'b011111001000;
        mem[5739] = 12'b011111000111;
        mem[5740] = 12'b011111000111;
        mem[5741] = 12'b011111000111;
        mem[5742] = 12'b011111000111;
        mem[5743] = 12'b011111000111;
        mem[5744] = 12'b011111000111;
        mem[5745] = 12'b011111000111;
        mem[5746] = 12'b011111000110;
        mem[5747] = 12'b011111000110;
        mem[5748] = 12'b011111000110;
        mem[5749] = 12'b011111000110;
        mem[5750] = 12'b011111000110;
        mem[5751] = 12'b011111000110;
        mem[5752] = 12'b011111000110;
        mem[5753] = 12'b011111000101;
        mem[5754] = 12'b011111000101;
        mem[5755] = 12'b011111000101;
        mem[5756] = 12'b011111000101;
        mem[5757] = 12'b011111000101;
        mem[5758] = 12'b011111000101;
        mem[5759] = 12'b011111000100;
        mem[5760] = 12'b011111000100;
        mem[5761] = 12'b011111000100;
        mem[5762] = 12'b011111000100;
        mem[5763] = 12'b011111000100;
        mem[5764] = 12'b011111000100;
        mem[5765] = 12'b011111000100;
        mem[5766] = 12'b011111000011;
        mem[5767] = 12'b011111000011;
        mem[5768] = 12'b011111000011;
        mem[5769] = 12'b011111000011;
        mem[5770] = 12'b011111000011;
        mem[5771] = 12'b011111000011;
        mem[5772] = 12'b011111000011;
        mem[5773] = 12'b011111000010;
        mem[5774] = 12'b011111000010;
        mem[5775] = 12'b011111000010;
        mem[5776] = 12'b011111000010;
        mem[5777] = 12'b011111000010;
        mem[5778] = 12'b011111000010;
        mem[5779] = 12'b011111000001;
        mem[5780] = 12'b011111000001;
        mem[5781] = 12'b011111000001;
        mem[5782] = 12'b011111000001;
        mem[5783] = 12'b011111000001;
        mem[5784] = 12'b011111000001;
        mem[5785] = 12'b011111000000;
        mem[5786] = 12'b011111000000;
        mem[5787] = 12'b011111000000;
        mem[5788] = 12'b011111000000;
        mem[5789] = 12'b011111000000;
        mem[5790] = 12'b011111000000;
        mem[5791] = 12'b011111000000;
        mem[5792] = 12'b011110111111;
        mem[5793] = 12'b011110111111;
        mem[5794] = 12'b011110111111;
        mem[5795] = 12'b011110111111;
        mem[5796] = 12'b011110111111;
        mem[5797] = 12'b011110111111;
        mem[5798] = 12'b011110111110;
        mem[5799] = 12'b011110111110;
        mem[5800] = 12'b011110111110;
        mem[5801] = 12'b011110111110;
        mem[5802] = 12'b011110111110;
        mem[5803] = 12'b011110111110;
        mem[5804] = 12'b011110111101;
        mem[5805] = 12'b011110111101;
        mem[5806] = 12'b011110111101;
        mem[5807] = 12'b011110111101;
        mem[5808] = 12'b011110111101;
        mem[5809] = 12'b011110111101;
        mem[5810] = 12'b011110111100;
        mem[5811] = 12'b011110111100;
        mem[5812] = 12'b011110111100;
        mem[5813] = 12'b011110111100;
        mem[5814] = 12'b011110111100;
        mem[5815] = 12'b011110111100;
        mem[5816] = 12'b011110111100;
        mem[5817] = 12'b011110111011;
        mem[5818] = 12'b011110111011;
        mem[5819] = 12'b011110111011;
        mem[5820] = 12'b011110111011;
        mem[5821] = 12'b011110111011;
        mem[5822] = 12'b011110111011;
        mem[5823] = 12'b011110111010;
        mem[5824] = 12'b011110111010;
        mem[5825] = 12'b011110111010;
        mem[5826] = 12'b011110111010;
        mem[5827] = 12'b011110111010;
        mem[5828] = 12'b011110111010;
        mem[5829] = 12'b011110111001;
        mem[5830] = 12'b011110111001;
        mem[5831] = 12'b011110111001;
        mem[5832] = 12'b011110111001;
        mem[5833] = 12'b011110111001;
        mem[5834] = 12'b011110111001;
        mem[5835] = 12'b011110111000;
        mem[5836] = 12'b011110111000;
        mem[5837] = 12'b011110111000;
        mem[5838] = 12'b011110111000;
        mem[5839] = 12'b011110111000;
        mem[5840] = 12'b011110111000;
        mem[5841] = 12'b011110110111;
        mem[5842] = 12'b011110110111;
        mem[5843] = 12'b011110110111;
        mem[5844] = 12'b011110110111;
        mem[5845] = 12'b011110110111;
        mem[5846] = 12'b011110110111;
        mem[5847] = 12'b011110110110;
        mem[5848] = 12'b011110110110;
        mem[5849] = 12'b011110110110;
        mem[5850] = 12'b011110110110;
        mem[5851] = 12'b011110110110;
        mem[5852] = 12'b011110110110;
        mem[5853] = 12'b011110110101;
        mem[5854] = 12'b011110110101;
        mem[5855] = 12'b011110110101;
        mem[5856] = 12'b011110110101;
        mem[5857] = 12'b011110110101;
        mem[5858] = 12'b011110110100;
        mem[5859] = 12'b011110110100;
        mem[5860] = 12'b011110110100;
        mem[5861] = 12'b011110110100;
        mem[5862] = 12'b011110110100;
        mem[5863] = 12'b011110110100;
        mem[5864] = 12'b011110110011;
        mem[5865] = 12'b011110110011;
        mem[5866] = 12'b011110110011;
        mem[5867] = 12'b011110110011;
        mem[5868] = 12'b011110110011;
        mem[5869] = 12'b011110110011;
        mem[5870] = 12'b011110110010;
        mem[5871] = 12'b011110110010;
        mem[5872] = 12'b011110110010;
        mem[5873] = 12'b011110110010;
        mem[5874] = 12'b011110110010;
        mem[5875] = 12'b011110110010;
        mem[5876] = 12'b011110110001;
        mem[5877] = 12'b011110110001;
        mem[5878] = 12'b011110110001;
        mem[5879] = 12'b011110110001;
        mem[5880] = 12'b011110110001;
        mem[5881] = 12'b011110110000;
        mem[5882] = 12'b011110110000;
        mem[5883] = 12'b011110110000;
        mem[5884] = 12'b011110110000;
        mem[5885] = 12'b011110110000;
        mem[5886] = 12'b011110110000;
        mem[5887] = 12'b011110101111;
        mem[5888] = 12'b011110101111;
        mem[5889] = 12'b011110101111;
        mem[5890] = 12'b011110101111;
        mem[5891] = 12'b011110101111;
        mem[5892] = 12'b011110101111;
        mem[5893] = 12'b011110101110;
        mem[5894] = 12'b011110101110;
        mem[5895] = 12'b011110101110;
        mem[5896] = 12'b011110101110;
        mem[5897] = 12'b011110101110;
        mem[5898] = 12'b011110101101;
        mem[5899] = 12'b011110101101;
        mem[5900] = 12'b011110101101;
        mem[5901] = 12'b011110101101;
        mem[5902] = 12'b011110101101;
        mem[5903] = 12'b011110101101;
        mem[5904] = 12'b011110101100;
        mem[5905] = 12'b011110101100;
        mem[5906] = 12'b011110101100;
        mem[5907] = 12'b011110101100;
        mem[5908] = 12'b011110101100;
        mem[5909] = 12'b011110101011;
        mem[5910] = 12'b011110101011;
        mem[5911] = 12'b011110101011;
        mem[5912] = 12'b011110101011;
        mem[5913] = 12'b011110101011;
        mem[5914] = 12'b011110101011;
        mem[5915] = 12'b011110101010;
        mem[5916] = 12'b011110101010;
        mem[5917] = 12'b011110101010;
        mem[5918] = 12'b011110101010;
        mem[5919] = 12'b011110101010;
        mem[5920] = 12'b011110101001;
        mem[5921] = 12'b011110101001;
        mem[5922] = 12'b011110101001;
        mem[5923] = 12'b011110101001;
        mem[5924] = 12'b011110101001;
        mem[5925] = 12'b011110101001;
        mem[5926] = 12'b011110101000;
        mem[5927] = 12'b011110101000;
        mem[5928] = 12'b011110101000;
        mem[5929] = 12'b011110101000;
        mem[5930] = 12'b011110101000;
        mem[5931] = 12'b011110100111;
        mem[5932] = 12'b011110100111;
        mem[5933] = 12'b011110100111;
        mem[5934] = 12'b011110100111;
        mem[5935] = 12'b011110100111;
        mem[5936] = 12'b011110100111;
        mem[5937] = 12'b011110100110;
        mem[5938] = 12'b011110100110;
        mem[5939] = 12'b011110100110;
        mem[5940] = 12'b011110100110;
        mem[5941] = 12'b011110100110;
        mem[5942] = 12'b011110100101;
        mem[5943] = 12'b011110100101;
        mem[5944] = 12'b011110100101;
        mem[5945] = 12'b011110100101;
        mem[5946] = 12'b011110100101;
        mem[5947] = 12'b011110100100;
        mem[5948] = 12'b011110100100;
        mem[5949] = 12'b011110100100;
        mem[5950] = 12'b011110100100;
        mem[5951] = 12'b011110100100;
        mem[5952] = 12'b011110100100;
        mem[5953] = 12'b011110100011;
        mem[5954] = 12'b011110100011;
        mem[5955] = 12'b011110100011;
        mem[5956] = 12'b011110100011;
        mem[5957] = 12'b011110100011;
        mem[5958] = 12'b011110100010;
        mem[5959] = 12'b011110100010;
        mem[5960] = 12'b011110100010;
        mem[5961] = 12'b011110100010;
        mem[5962] = 12'b011110100010;
        mem[5963] = 12'b011110100001;
        mem[5964] = 12'b011110100001;
        mem[5965] = 12'b011110100001;
        mem[5966] = 12'b011110100001;
        mem[5967] = 12'b011110100001;
        mem[5968] = 12'b011110100000;
        mem[5969] = 12'b011110100000;
        mem[5970] = 12'b011110100000;
        mem[5971] = 12'b011110100000;
        mem[5972] = 12'b011110100000;
        mem[5973] = 12'b011110011111;
        mem[5974] = 12'b011110011111;
        mem[5975] = 12'b011110011111;
        mem[5976] = 12'b011110011111;
        mem[5977] = 12'b011110011111;
        mem[5978] = 12'b011110011111;
        mem[5979] = 12'b011110011110;
        mem[5980] = 12'b011110011110;
        mem[5981] = 12'b011110011110;
        mem[5982] = 12'b011110011110;
        mem[5983] = 12'b011110011110;
        mem[5984] = 12'b011110011101;
        mem[5985] = 12'b011110011101;
        mem[5986] = 12'b011110011101;
        mem[5987] = 12'b011110011101;
        mem[5988] = 12'b011110011101;
        mem[5989] = 12'b011110011100;
        mem[5990] = 12'b011110011100;
        mem[5991] = 12'b011110011100;
        mem[5992] = 12'b011110011100;
        mem[5993] = 12'b011110011100;
        mem[5994] = 12'b011110011011;
        mem[5995] = 12'b011110011011;
        mem[5996] = 12'b011110011011;
        mem[5997] = 12'b011110011011;
        mem[5998] = 12'b011110011011;
        mem[5999] = 12'b011110011010;
        mem[6000] = 12'b011110011010;
        mem[6001] = 12'b011110011010;
        mem[6002] = 12'b011110011010;
        mem[6003] = 12'b011110011010;
        mem[6004] = 12'b011110011001;
        mem[6005] = 12'b011110011001;
        mem[6006] = 12'b011110011001;
        mem[6007] = 12'b011110011001;
        mem[6008] = 12'b011110011001;
        mem[6009] = 12'b011110011000;
        mem[6010] = 12'b011110011000;
        mem[6011] = 12'b011110011000;
        mem[6012] = 12'b011110011000;
        mem[6013] = 12'b011110011000;
        mem[6014] = 12'b011110010111;
        mem[6015] = 12'b011110010111;
        mem[6016] = 12'b011110010111;
        mem[6017] = 12'b011110010111;
        mem[6018] = 12'b011110010111;
        mem[6019] = 12'b011110010110;
        mem[6020] = 12'b011110010110;
        mem[6021] = 12'b011110010110;
        mem[6022] = 12'b011110010110;
        mem[6023] = 12'b011110010110;
        mem[6024] = 12'b011110010101;
        mem[6025] = 12'b011110010101;
        mem[6026] = 12'b011110010101;
        mem[6027] = 12'b011110010101;
        mem[6028] = 12'b011110010101;
        mem[6029] = 12'b011110010100;
        mem[6030] = 12'b011110010100;
        mem[6031] = 12'b011110010100;
        mem[6032] = 12'b011110010100;
        mem[6033] = 12'b011110010100;
        mem[6034] = 12'b011110010011;
        mem[6035] = 12'b011110010011;
        mem[6036] = 12'b011110010011;
        mem[6037] = 12'b011110010011;
        mem[6038] = 12'b011110010010;
        mem[6039] = 12'b011110010010;
        mem[6040] = 12'b011110010010;
        mem[6041] = 12'b011110010010;
        mem[6042] = 12'b011110010010;
        mem[6043] = 12'b011110010001;
        mem[6044] = 12'b011110010001;
        mem[6045] = 12'b011110010001;
        mem[6046] = 12'b011110010001;
        mem[6047] = 12'b011110010001;
        mem[6048] = 12'b011110010000;
        mem[6049] = 12'b011110010000;
        mem[6050] = 12'b011110010000;
        mem[6051] = 12'b011110010000;
        mem[6052] = 12'b011110010000;
        mem[6053] = 12'b011110001111;
        mem[6054] = 12'b011110001111;
        mem[6055] = 12'b011110001111;
        mem[6056] = 12'b011110001111;
        mem[6057] = 12'b011110001111;
        mem[6058] = 12'b011110001110;
        mem[6059] = 12'b011110001110;
        mem[6060] = 12'b011110001110;
        mem[6061] = 12'b011110001110;
        mem[6062] = 12'b011110001101;
        mem[6063] = 12'b011110001101;
        mem[6064] = 12'b011110001101;
        mem[6065] = 12'b011110001101;
        mem[6066] = 12'b011110001101;
        mem[6067] = 12'b011110001100;
        mem[6068] = 12'b011110001100;
        mem[6069] = 12'b011110001100;
        mem[6070] = 12'b011110001100;
        mem[6071] = 12'b011110001100;
        mem[6072] = 12'b011110001011;
        mem[6073] = 12'b011110001011;
        mem[6074] = 12'b011110001011;
        mem[6075] = 12'b011110001011;
        mem[6076] = 12'b011110001011;
        mem[6077] = 12'b011110001010;
        mem[6078] = 12'b011110001010;
        mem[6079] = 12'b011110001010;
        mem[6080] = 12'b011110001010;
        mem[6081] = 12'b011110001001;
        mem[6082] = 12'b011110001001;
        mem[6083] = 12'b011110001001;
        mem[6084] = 12'b011110001001;
        mem[6085] = 12'b011110001001;
        mem[6086] = 12'b011110001000;
        mem[6087] = 12'b011110001000;
        mem[6088] = 12'b011110001000;
        mem[6089] = 12'b011110001000;
        mem[6090] = 12'b011110001000;
        mem[6091] = 12'b011110000111;
        mem[6092] = 12'b011110000111;
        mem[6093] = 12'b011110000111;
        mem[6094] = 12'b011110000111;
        mem[6095] = 12'b011110000110;
        mem[6096] = 12'b011110000110;
        mem[6097] = 12'b011110000110;
        mem[6098] = 12'b011110000110;
        mem[6099] = 12'b011110000110;
        mem[6100] = 12'b011110000101;
        mem[6101] = 12'b011110000101;
        mem[6102] = 12'b011110000101;
        mem[6103] = 12'b011110000101;
        mem[6104] = 12'b011110000100;
        mem[6105] = 12'b011110000100;
        mem[6106] = 12'b011110000100;
        mem[6107] = 12'b011110000100;
        mem[6108] = 12'b011110000100;
        mem[6109] = 12'b011110000011;
        mem[6110] = 12'b011110000011;
        mem[6111] = 12'b011110000011;
        mem[6112] = 12'b011110000011;
        mem[6113] = 12'b011110000011;
        mem[6114] = 12'b011110000010;
        mem[6115] = 12'b011110000010;
        mem[6116] = 12'b011110000010;
        mem[6117] = 12'b011110000010;
        mem[6118] = 12'b011110000001;
        mem[6119] = 12'b011110000001;
        mem[6120] = 12'b011110000001;
        mem[6121] = 12'b011110000001;
        mem[6122] = 12'b011110000001;
        mem[6123] = 12'b011110000000;
        mem[6124] = 12'b011110000000;
        mem[6125] = 12'b011110000000;
        mem[6126] = 12'b011110000000;
        mem[6127] = 12'b011101111111;
        mem[6128] = 12'b011101111111;
        mem[6129] = 12'b011101111111;
        mem[6130] = 12'b011101111111;
        mem[6131] = 12'b011101111111;
        mem[6132] = 12'b011101111110;
        mem[6133] = 12'b011101111110;
        mem[6134] = 12'b011101111110;
        mem[6135] = 12'b011101111110;
        mem[6136] = 12'b011101111101;
        mem[6137] = 12'b011101111101;
        mem[6138] = 12'b011101111101;
        mem[6139] = 12'b011101111101;
        mem[6140] = 12'b011101111100;
        mem[6141] = 12'b011101111100;
        mem[6142] = 12'b011101111100;
        mem[6143] = 12'b011101111100;
        mem[6144] = 12'b011101111100;
        mem[6145] = 12'b011101111011;
        mem[6146] = 12'b011101111011;
        mem[6147] = 12'b011101111011;
        mem[6148] = 12'b011101111011;
        mem[6149] = 12'b011101111010;
        mem[6150] = 12'b011101111010;
        mem[6151] = 12'b011101111010;
        mem[6152] = 12'b011101111010;
        mem[6153] = 12'b011101111010;
        mem[6154] = 12'b011101111001;
        mem[6155] = 12'b011101111001;
        mem[6156] = 12'b011101111001;
        mem[6157] = 12'b011101111001;
        mem[6158] = 12'b011101111000;
        mem[6159] = 12'b011101111000;
        mem[6160] = 12'b011101111000;
        mem[6161] = 12'b011101111000;
        mem[6162] = 12'b011101110111;
        mem[6163] = 12'b011101110111;
        mem[6164] = 12'b011101110111;
        mem[6165] = 12'b011101110111;
        mem[6166] = 12'b011101110111;
        mem[6167] = 12'b011101110110;
        mem[6168] = 12'b011101110110;
        mem[6169] = 12'b011101110110;
        mem[6170] = 12'b011101110110;
        mem[6171] = 12'b011101110101;
        mem[6172] = 12'b011101110101;
        mem[6173] = 12'b011101110101;
        mem[6174] = 12'b011101110101;
        mem[6175] = 12'b011101110100;
        mem[6176] = 12'b011101110100;
        mem[6177] = 12'b011101110100;
        mem[6178] = 12'b011101110100;
        mem[6179] = 12'b011101110100;
        mem[6180] = 12'b011101110011;
        mem[6181] = 12'b011101110011;
        mem[6182] = 12'b011101110011;
        mem[6183] = 12'b011101110011;
        mem[6184] = 12'b011101110010;
        mem[6185] = 12'b011101110010;
        mem[6186] = 12'b011101110010;
        mem[6187] = 12'b011101110010;
        mem[6188] = 12'b011101110001;
        mem[6189] = 12'b011101110001;
        mem[6190] = 12'b011101110001;
        mem[6191] = 12'b011101110001;
        mem[6192] = 12'b011101110000;
        mem[6193] = 12'b011101110000;
        mem[6194] = 12'b011101110000;
        mem[6195] = 12'b011101110000;
        mem[6196] = 12'b011101110000;
        mem[6197] = 12'b011101101111;
        mem[6198] = 12'b011101101111;
        mem[6199] = 12'b011101101111;
        mem[6200] = 12'b011101101111;
        mem[6201] = 12'b011101101110;
        mem[6202] = 12'b011101101110;
        mem[6203] = 12'b011101101110;
        mem[6204] = 12'b011101101110;
        mem[6205] = 12'b011101101101;
        mem[6206] = 12'b011101101101;
        mem[6207] = 12'b011101101101;
        mem[6208] = 12'b011101101101;
        mem[6209] = 12'b011101101100;
        mem[6210] = 12'b011101101100;
        mem[6211] = 12'b011101101100;
        mem[6212] = 12'b011101101100;
        mem[6213] = 12'b011101101100;
        mem[6214] = 12'b011101101011;
        mem[6215] = 12'b011101101011;
        mem[6216] = 12'b011101101011;
        mem[6217] = 12'b011101101011;
        mem[6218] = 12'b011101101010;
        mem[6219] = 12'b011101101010;
        mem[6220] = 12'b011101101010;
        mem[6221] = 12'b011101101010;
        mem[6222] = 12'b011101101001;
        mem[6223] = 12'b011101101001;
        mem[6224] = 12'b011101101001;
        mem[6225] = 12'b011101101001;
        mem[6226] = 12'b011101101000;
        mem[6227] = 12'b011101101000;
        mem[6228] = 12'b011101101000;
        mem[6229] = 12'b011101101000;
        mem[6230] = 12'b011101100111;
        mem[6231] = 12'b011101100111;
        mem[6232] = 12'b011101100111;
        mem[6233] = 12'b011101100111;
        mem[6234] = 12'b011101100110;
        mem[6235] = 12'b011101100110;
        mem[6236] = 12'b011101100110;
        mem[6237] = 12'b011101100110;
        mem[6238] = 12'b011101100101;
        mem[6239] = 12'b011101100101;
        mem[6240] = 12'b011101100101;
        mem[6241] = 12'b011101100101;
        mem[6242] = 12'b011101100100;
        mem[6243] = 12'b011101100100;
        mem[6244] = 12'b011101100100;
        mem[6245] = 12'b011101100100;
        mem[6246] = 12'b011101100100;
        mem[6247] = 12'b011101100011;
        mem[6248] = 12'b011101100011;
        mem[6249] = 12'b011101100011;
        mem[6250] = 12'b011101100011;
        mem[6251] = 12'b011101100010;
        mem[6252] = 12'b011101100010;
        mem[6253] = 12'b011101100010;
        mem[6254] = 12'b011101100010;
        mem[6255] = 12'b011101100001;
        mem[6256] = 12'b011101100001;
        mem[6257] = 12'b011101100001;
        mem[6258] = 12'b011101100001;
        mem[6259] = 12'b011101100000;
        mem[6260] = 12'b011101100000;
        mem[6261] = 12'b011101100000;
        mem[6262] = 12'b011101100000;
        mem[6263] = 12'b011101011111;
        mem[6264] = 12'b011101011111;
        mem[6265] = 12'b011101011111;
        mem[6266] = 12'b011101011111;
        mem[6267] = 12'b011101011110;
        mem[6268] = 12'b011101011110;
        mem[6269] = 12'b011101011110;
        mem[6270] = 12'b011101011110;
        mem[6271] = 12'b011101011101;
        mem[6272] = 12'b011101011101;
        mem[6273] = 12'b011101011101;
        mem[6274] = 12'b011101011101;
        mem[6275] = 12'b011101011100;
        mem[6276] = 12'b011101011100;
        mem[6277] = 12'b011101011100;
        mem[6278] = 12'b011101011100;
        mem[6279] = 12'b011101011011;
        mem[6280] = 12'b011101011011;
        mem[6281] = 12'b011101011011;
        mem[6282] = 12'b011101011011;
        mem[6283] = 12'b011101011010;
        mem[6284] = 12'b011101011010;
        mem[6285] = 12'b011101011010;
        mem[6286] = 12'b011101011010;
        mem[6287] = 12'b011101011001;
        mem[6288] = 12'b011101011001;
        mem[6289] = 12'b011101011001;
        mem[6290] = 12'b011101011001;
        mem[6291] = 12'b011101011000;
        mem[6292] = 12'b011101011000;
        mem[6293] = 12'b011101011000;
        mem[6294] = 12'b011101011000;
        mem[6295] = 12'b011101010111;
        mem[6296] = 12'b011101010111;
        mem[6297] = 12'b011101010111;
        mem[6298] = 12'b011101010110;
        mem[6299] = 12'b011101010110;
        mem[6300] = 12'b011101010110;
        mem[6301] = 12'b011101010110;
        mem[6302] = 12'b011101010101;
        mem[6303] = 12'b011101010101;
        mem[6304] = 12'b011101010101;
        mem[6305] = 12'b011101010101;
        mem[6306] = 12'b011101010100;
        mem[6307] = 12'b011101010100;
        mem[6308] = 12'b011101010100;
        mem[6309] = 12'b011101010100;
        mem[6310] = 12'b011101010011;
        mem[6311] = 12'b011101010011;
        mem[6312] = 12'b011101010011;
        mem[6313] = 12'b011101010011;
        mem[6314] = 12'b011101010010;
        mem[6315] = 12'b011101010010;
        mem[6316] = 12'b011101010010;
        mem[6317] = 12'b011101010010;
        mem[6318] = 12'b011101010001;
        mem[6319] = 12'b011101010001;
        mem[6320] = 12'b011101010001;
        mem[6321] = 12'b011101010001;
        mem[6322] = 12'b011101010000;
        mem[6323] = 12'b011101010000;
        mem[6324] = 12'b011101010000;
        mem[6325] = 12'b011101010000;
        mem[6326] = 12'b011101001111;
        mem[6327] = 12'b011101001111;
        mem[6328] = 12'b011101001111;
        mem[6329] = 12'b011101001110;
        mem[6330] = 12'b011101001110;
        mem[6331] = 12'b011101001110;
        mem[6332] = 12'b011101001110;
        mem[6333] = 12'b011101001101;
        mem[6334] = 12'b011101001101;
        mem[6335] = 12'b011101001101;
        mem[6336] = 12'b011101001101;
        mem[6337] = 12'b011101001100;
        mem[6338] = 12'b011101001100;
        mem[6339] = 12'b011101001100;
        mem[6340] = 12'b011101001100;
        mem[6341] = 12'b011101001011;
        mem[6342] = 12'b011101001011;
        mem[6343] = 12'b011101001011;
        mem[6344] = 12'b011101001011;
        mem[6345] = 12'b011101001010;
        mem[6346] = 12'b011101001010;
        mem[6347] = 12'b011101001010;
        mem[6348] = 12'b011101001010;
        mem[6349] = 12'b011101001001;
        mem[6350] = 12'b011101001001;
        mem[6351] = 12'b011101001001;
        mem[6352] = 12'b011101001000;
        mem[6353] = 12'b011101001000;
        mem[6354] = 12'b011101001000;
        mem[6355] = 12'b011101001000;
        mem[6356] = 12'b011101000111;
        mem[6357] = 12'b011101000111;
        mem[6358] = 12'b011101000111;
        mem[6359] = 12'b011101000111;
        mem[6360] = 12'b011101000110;
        mem[6361] = 12'b011101000110;
        mem[6362] = 12'b011101000110;
        mem[6363] = 12'b011101000110;
        mem[6364] = 12'b011101000101;
        mem[6365] = 12'b011101000101;
        mem[6366] = 12'b011101000101;
        mem[6367] = 12'b011101000100;
        mem[6368] = 12'b011101000100;
        mem[6369] = 12'b011101000100;
        mem[6370] = 12'b011101000100;
        mem[6371] = 12'b011101000011;
        mem[6372] = 12'b011101000011;
        mem[6373] = 12'b011101000011;
        mem[6374] = 12'b011101000011;
        mem[6375] = 12'b011101000010;
        mem[6376] = 12'b011101000010;
        mem[6377] = 12'b011101000010;
        mem[6378] = 12'b011101000001;
        mem[6379] = 12'b011101000001;
        mem[6380] = 12'b011101000001;
        mem[6381] = 12'b011101000001;
        mem[6382] = 12'b011101000000;
        mem[6383] = 12'b011101000000;
        mem[6384] = 12'b011101000000;
        mem[6385] = 12'b011101000000;
        mem[6386] = 12'b011100111111;
        mem[6387] = 12'b011100111111;
        mem[6388] = 12'b011100111111;
        mem[6389] = 12'b011100111111;
        mem[6390] = 12'b011100111110;
        mem[6391] = 12'b011100111110;
        mem[6392] = 12'b011100111110;
        mem[6393] = 12'b011100111101;
        mem[6394] = 12'b011100111101;
        mem[6395] = 12'b011100111101;
        mem[6396] = 12'b011100111101;
        mem[6397] = 12'b011100111100;
        mem[6398] = 12'b011100111100;
        mem[6399] = 12'b011100111100;
        mem[6400] = 12'b011100111100;
        mem[6401] = 12'b011100111011;
        mem[6402] = 12'b011100111011;
        mem[6403] = 12'b011100111011;
        mem[6404] = 12'b011100111010;
        mem[6405] = 12'b011100111010;
        mem[6406] = 12'b011100111010;
        mem[6407] = 12'b011100111010;
        mem[6408] = 12'b011100111001;
        mem[6409] = 12'b011100111001;
        mem[6410] = 12'b011100111001;
        mem[6411] = 12'b011100111000;
        mem[6412] = 12'b011100111000;
        mem[6413] = 12'b011100111000;
        mem[6414] = 12'b011100111000;
        mem[6415] = 12'b011100110111;
        mem[6416] = 12'b011100110111;
        mem[6417] = 12'b011100110111;
        mem[6418] = 12'b011100110111;
        mem[6419] = 12'b011100110110;
        mem[6420] = 12'b011100110110;
        mem[6421] = 12'b011100110110;
        mem[6422] = 12'b011100110101;
        mem[6423] = 12'b011100110101;
        mem[6424] = 12'b011100110101;
        mem[6425] = 12'b011100110101;
        mem[6426] = 12'b011100110100;
        mem[6427] = 12'b011100110100;
        mem[6428] = 12'b011100110100;
        mem[6429] = 12'b011100110011;
        mem[6430] = 12'b011100110011;
        mem[6431] = 12'b011100110011;
        mem[6432] = 12'b011100110011;
        mem[6433] = 12'b011100110010;
        mem[6434] = 12'b011100110010;
        mem[6435] = 12'b011100110010;
        mem[6436] = 12'b011100110010;
        mem[6437] = 12'b011100110001;
        mem[6438] = 12'b011100110001;
        mem[6439] = 12'b011100110001;
        mem[6440] = 12'b011100110000;
        mem[6441] = 12'b011100110000;
        mem[6442] = 12'b011100110000;
        mem[6443] = 12'b011100110000;
        mem[6444] = 12'b011100101111;
        mem[6445] = 12'b011100101111;
        mem[6446] = 12'b011100101111;
        mem[6447] = 12'b011100101110;
        mem[6448] = 12'b011100101110;
        mem[6449] = 12'b011100101110;
        mem[6450] = 12'b011100101110;
        mem[6451] = 12'b011100101101;
        mem[6452] = 12'b011100101101;
        mem[6453] = 12'b011100101101;
        mem[6454] = 12'b011100101100;
        mem[6455] = 12'b011100101100;
        mem[6456] = 12'b011100101100;
        mem[6457] = 12'b011100101100;
        mem[6458] = 12'b011100101011;
        mem[6459] = 12'b011100101011;
        mem[6460] = 12'b011100101011;
        mem[6461] = 12'b011100101010;
        mem[6462] = 12'b011100101010;
        mem[6463] = 12'b011100101010;
        mem[6464] = 12'b011100101010;
        mem[6465] = 12'b011100101001;
        mem[6466] = 12'b011100101001;
        mem[6467] = 12'b011100101001;
        mem[6468] = 12'b011100101000;
        mem[6469] = 12'b011100101000;
        mem[6470] = 12'b011100101000;
        mem[6471] = 12'b011100101000;
        mem[6472] = 12'b011100100111;
        mem[6473] = 12'b011100100111;
        mem[6474] = 12'b011100100111;
        mem[6475] = 12'b011100100110;
        mem[6476] = 12'b011100100110;
        mem[6477] = 12'b011100100110;
        mem[6478] = 12'b011100100110;
        mem[6479] = 12'b011100100101;
        mem[6480] = 12'b011100100101;
        mem[6481] = 12'b011100100101;
        mem[6482] = 12'b011100100100;
        mem[6483] = 12'b011100100100;
        mem[6484] = 12'b011100100100;
        mem[6485] = 12'b011100100100;
        mem[6486] = 12'b011100100011;
        mem[6487] = 12'b011100100011;
        mem[6488] = 12'b011100100011;
        mem[6489] = 12'b011100100010;
        mem[6490] = 12'b011100100010;
        mem[6491] = 12'b011100100010;
        mem[6492] = 12'b011100100010;
        mem[6493] = 12'b011100100001;
        mem[6494] = 12'b011100100001;
        mem[6495] = 12'b011100100001;
        mem[6496] = 12'b011100100000;
        mem[6497] = 12'b011100100000;
        mem[6498] = 12'b011100100000;
        mem[6499] = 12'b011100011111;
        mem[6500] = 12'b011100011111;
        mem[6501] = 12'b011100011111;
        mem[6502] = 12'b011100011111;
        mem[6503] = 12'b011100011110;
        mem[6504] = 12'b011100011110;
        mem[6505] = 12'b011100011110;
        mem[6506] = 12'b011100011101;
        mem[6507] = 12'b011100011101;
        mem[6508] = 12'b011100011101;
        mem[6509] = 12'b011100011101;
        mem[6510] = 12'b011100011100;
        mem[6511] = 12'b011100011100;
        mem[6512] = 12'b011100011100;
        mem[6513] = 12'b011100011011;
        mem[6514] = 12'b011100011011;
        mem[6515] = 12'b011100011011;
        mem[6516] = 12'b011100011011;
        mem[6517] = 12'b011100011010;
        mem[6518] = 12'b011100011010;
        mem[6519] = 12'b011100011010;
        mem[6520] = 12'b011100011001;
        mem[6521] = 12'b011100011001;
        mem[6522] = 12'b011100011001;
        mem[6523] = 12'b011100011000;
        mem[6524] = 12'b011100011000;
        mem[6525] = 12'b011100011000;
        mem[6526] = 12'b011100011000;
        mem[6527] = 12'b011100010111;
        mem[6528] = 12'b011100010111;
        mem[6529] = 12'b011100010111;
        mem[6530] = 12'b011100010110;
        mem[6531] = 12'b011100010110;
        mem[6532] = 12'b011100010110;
        mem[6533] = 12'b011100010101;
        mem[6534] = 12'b011100010101;
        mem[6535] = 12'b011100010101;
        mem[6536] = 12'b011100010101;
        mem[6537] = 12'b011100010100;
        mem[6538] = 12'b011100010100;
        mem[6539] = 12'b011100010100;
        mem[6540] = 12'b011100010011;
        mem[6541] = 12'b011100010011;
        mem[6542] = 12'b011100010011;
        mem[6543] = 12'b011100010010;
        mem[6544] = 12'b011100010010;
        mem[6545] = 12'b011100010010;
        mem[6546] = 12'b011100010010;
        mem[6547] = 12'b011100010001;
        mem[6548] = 12'b011100010001;
        mem[6549] = 12'b011100010001;
        mem[6550] = 12'b011100010000;
        mem[6551] = 12'b011100010000;
        mem[6552] = 12'b011100010000;
        mem[6553] = 12'b011100001111;
        mem[6554] = 12'b011100001111;
        mem[6555] = 12'b011100001111;
        mem[6556] = 12'b011100001111;
        mem[6557] = 12'b011100001110;
        mem[6558] = 12'b011100001110;
        mem[6559] = 12'b011100001110;
        mem[6560] = 12'b011100001101;
        mem[6561] = 12'b011100001101;
        mem[6562] = 12'b011100001101;
        mem[6563] = 12'b011100001100;
        mem[6564] = 12'b011100001100;
        mem[6565] = 12'b011100001100;
        mem[6566] = 12'b011100001100;
        mem[6567] = 12'b011100001011;
        mem[6568] = 12'b011100001011;
        mem[6569] = 12'b011100001011;
        mem[6570] = 12'b011100001010;
        mem[6571] = 12'b011100001010;
        mem[6572] = 12'b011100001010;
        mem[6573] = 12'b011100001001;
        mem[6574] = 12'b011100001001;
        mem[6575] = 12'b011100001001;
        mem[6576] = 12'b011100001000;
        mem[6577] = 12'b011100001000;
        mem[6578] = 12'b011100001000;
        mem[6579] = 12'b011100001000;
        mem[6580] = 12'b011100000111;
        mem[6581] = 12'b011100000111;
        mem[6582] = 12'b011100000111;
        mem[6583] = 12'b011100000110;
        mem[6584] = 12'b011100000110;
        mem[6585] = 12'b011100000110;
        mem[6586] = 12'b011100000101;
        mem[6587] = 12'b011100000101;
        mem[6588] = 12'b011100000101;
        mem[6589] = 12'b011100000100;
        mem[6590] = 12'b011100000100;
        mem[6591] = 12'b011100000100;
        mem[6592] = 12'b011100000100;
        mem[6593] = 12'b011100000011;
        mem[6594] = 12'b011100000011;
        mem[6595] = 12'b011100000011;
        mem[6596] = 12'b011100000010;
        mem[6597] = 12'b011100000010;
        mem[6598] = 12'b011100000010;
        mem[6599] = 12'b011100000001;
        mem[6600] = 12'b011100000001;
        mem[6601] = 12'b011100000001;
        mem[6602] = 12'b011100000000;
        mem[6603] = 12'b011100000000;
        mem[6604] = 12'b011100000000;
        mem[6605] = 12'b011100000000;
        mem[6606] = 12'b011011111111;
        mem[6607] = 12'b011011111111;
        mem[6608] = 12'b011011111111;
        mem[6609] = 12'b011011111110;
        mem[6610] = 12'b011011111110;
        mem[6611] = 12'b011011111110;
        mem[6612] = 12'b011011111101;
        mem[6613] = 12'b011011111101;
        mem[6614] = 12'b011011111101;
        mem[6615] = 12'b011011111100;
        mem[6616] = 12'b011011111100;
        mem[6617] = 12'b011011111100;
        mem[6618] = 12'b011011111011;
        mem[6619] = 12'b011011111011;
        mem[6620] = 12'b011011111011;
        mem[6621] = 12'b011011111011;
        mem[6622] = 12'b011011111010;
        mem[6623] = 12'b011011111010;
        mem[6624] = 12'b011011111010;
        mem[6625] = 12'b011011111001;
        mem[6626] = 12'b011011111001;
        mem[6627] = 12'b011011111001;
        mem[6628] = 12'b011011111000;
        mem[6629] = 12'b011011111000;
        mem[6630] = 12'b011011111000;
        mem[6631] = 12'b011011110111;
        mem[6632] = 12'b011011110111;
        mem[6633] = 12'b011011110111;
        mem[6634] = 12'b011011110110;
        mem[6635] = 12'b011011110110;
        mem[6636] = 12'b011011110110;
        mem[6637] = 12'b011011110110;
        mem[6638] = 12'b011011110101;
        mem[6639] = 12'b011011110101;
        mem[6640] = 12'b011011110101;
        mem[6641] = 12'b011011110100;
        mem[6642] = 12'b011011110100;
        mem[6643] = 12'b011011110100;
        mem[6644] = 12'b011011110011;
        mem[6645] = 12'b011011110011;
        mem[6646] = 12'b011011110011;
        mem[6647] = 12'b011011110010;
        mem[6648] = 12'b011011110010;
        mem[6649] = 12'b011011110010;
        mem[6650] = 12'b011011110001;
        mem[6651] = 12'b011011110001;
        mem[6652] = 12'b011011110001;
        mem[6653] = 12'b011011110000;
        mem[6654] = 12'b011011110000;
        mem[6655] = 12'b011011110000;
        mem[6656] = 12'b011011101111;
        mem[6657] = 12'b011011101111;
        mem[6658] = 12'b011011101111;
        mem[6659] = 12'b011011101111;
        mem[6660] = 12'b011011101110;
        mem[6661] = 12'b011011101110;
        mem[6662] = 12'b011011101110;
        mem[6663] = 12'b011011101101;
        mem[6664] = 12'b011011101101;
        mem[6665] = 12'b011011101101;
        mem[6666] = 12'b011011101100;
        mem[6667] = 12'b011011101100;
        mem[6668] = 12'b011011101100;
        mem[6669] = 12'b011011101011;
        mem[6670] = 12'b011011101011;
        mem[6671] = 12'b011011101011;
        mem[6672] = 12'b011011101010;
        mem[6673] = 12'b011011101010;
        mem[6674] = 12'b011011101010;
        mem[6675] = 12'b011011101001;
        mem[6676] = 12'b011011101001;
        mem[6677] = 12'b011011101001;
        mem[6678] = 12'b011011101000;
        mem[6679] = 12'b011011101000;
        mem[6680] = 12'b011011101000;
        mem[6681] = 12'b011011100111;
        mem[6682] = 12'b011011100111;
        mem[6683] = 12'b011011100111;
        mem[6684] = 12'b011011100110;
        mem[6685] = 12'b011011100110;
        mem[6686] = 12'b011011100110;
        mem[6687] = 12'b011011100101;
        mem[6688] = 12'b011011100101;
        mem[6689] = 12'b011011100101;
        mem[6690] = 12'b011011100100;
        mem[6691] = 12'b011011100100;
        mem[6692] = 12'b011011100100;
        mem[6693] = 12'b011011100100;
        mem[6694] = 12'b011011100011;
        mem[6695] = 12'b011011100011;
        mem[6696] = 12'b011011100011;
        mem[6697] = 12'b011011100010;
        mem[6698] = 12'b011011100010;
        mem[6699] = 12'b011011100010;
        mem[6700] = 12'b011011100001;
        mem[6701] = 12'b011011100001;
        mem[6702] = 12'b011011100001;
        mem[6703] = 12'b011011100000;
        mem[6704] = 12'b011011100000;
        mem[6705] = 12'b011011100000;
        mem[6706] = 12'b011011011111;
        mem[6707] = 12'b011011011111;
        mem[6708] = 12'b011011011111;
        mem[6709] = 12'b011011011110;
        mem[6710] = 12'b011011011110;
        mem[6711] = 12'b011011011110;
        mem[6712] = 12'b011011011101;
        mem[6713] = 12'b011011011101;
        mem[6714] = 12'b011011011101;
        mem[6715] = 12'b011011011100;
        mem[6716] = 12'b011011011100;
        mem[6717] = 12'b011011011100;
        mem[6718] = 12'b011011011011;
        mem[6719] = 12'b011011011011;
        mem[6720] = 12'b011011011011;
        mem[6721] = 12'b011011011010;
        mem[6722] = 12'b011011011010;
        mem[6723] = 12'b011011011010;
        mem[6724] = 12'b011011011001;
        mem[6725] = 12'b011011011001;
        mem[6726] = 12'b011011011001;
        mem[6727] = 12'b011011011000;
        mem[6728] = 12'b011011011000;
        mem[6729] = 12'b011011011000;
        mem[6730] = 12'b011011010111;
        mem[6731] = 12'b011011010111;
        mem[6732] = 12'b011011010111;
        mem[6733] = 12'b011011010110;
        mem[6734] = 12'b011011010110;
        mem[6735] = 12'b011011010110;
        mem[6736] = 12'b011011010101;
        mem[6737] = 12'b011011010101;
        mem[6738] = 12'b011011010101;
        mem[6739] = 12'b011011010100;
        mem[6740] = 12'b011011010100;
        mem[6741] = 12'b011011010100;
        mem[6742] = 12'b011011010011;
        mem[6743] = 12'b011011010011;
        mem[6744] = 12'b011011010011;
        mem[6745] = 12'b011011010010;
        mem[6746] = 12'b011011010010;
        mem[6747] = 12'b011011010010;
        mem[6748] = 12'b011011010001;
        mem[6749] = 12'b011011010001;
        mem[6750] = 12'b011011010001;
        mem[6751] = 12'b011011010000;
        mem[6752] = 12'b011011010000;
        mem[6753] = 12'b011011010000;
        mem[6754] = 12'b011011001111;
        mem[6755] = 12'b011011001111;
        mem[6756] = 12'b011011001111;
        mem[6757] = 12'b011011001110;
        mem[6758] = 12'b011011001110;
        mem[6759] = 12'b011011001110;
        mem[6760] = 12'b011011001101;
        mem[6761] = 12'b011011001101;
        mem[6762] = 12'b011011001101;
        mem[6763] = 12'b011011001100;
        mem[6764] = 12'b011011001100;
        mem[6765] = 12'b011011001100;
        mem[6766] = 12'b011011001011;
        mem[6767] = 12'b011011001011;
        mem[6768] = 12'b011011001011;
        mem[6769] = 12'b011011001010;
        mem[6770] = 12'b011011001010;
        mem[6771] = 12'b011011001010;
        mem[6772] = 12'b011011001001;
        mem[6773] = 12'b011011001001;
        mem[6774] = 12'b011011001001;
        mem[6775] = 12'b011011001000;
        mem[6776] = 12'b011011001000;
        mem[6777] = 12'b011011000111;
        mem[6778] = 12'b011011000111;
        mem[6779] = 12'b011011000111;
        mem[6780] = 12'b011011000110;
        mem[6781] = 12'b011011000110;
        mem[6782] = 12'b011011000110;
        mem[6783] = 12'b011011000101;
        mem[6784] = 12'b011011000101;
        mem[6785] = 12'b011011000101;
        mem[6786] = 12'b011011000100;
        mem[6787] = 12'b011011000100;
        mem[6788] = 12'b011011000100;
        mem[6789] = 12'b011011000011;
        mem[6790] = 12'b011011000011;
        mem[6791] = 12'b011011000011;
        mem[6792] = 12'b011011000010;
        mem[6793] = 12'b011011000010;
        mem[6794] = 12'b011011000010;
        mem[6795] = 12'b011011000001;
        mem[6796] = 12'b011011000001;
        mem[6797] = 12'b011011000001;
        mem[6798] = 12'b011011000000;
        mem[6799] = 12'b011011000000;
        mem[6800] = 12'b011011000000;
        mem[6801] = 12'b011010111111;
        mem[6802] = 12'b011010111111;
        mem[6803] = 12'b011010111111;
        mem[6804] = 12'b011010111110;
        mem[6805] = 12'b011010111110;
        mem[6806] = 12'b011010111110;
        mem[6807] = 12'b011010111101;
        mem[6808] = 12'b011010111101;
        mem[6809] = 12'b011010111100;
        mem[6810] = 12'b011010111100;
        mem[6811] = 12'b011010111100;
        mem[6812] = 12'b011010111011;
        mem[6813] = 12'b011010111011;
        mem[6814] = 12'b011010111011;
        mem[6815] = 12'b011010111010;
        mem[6816] = 12'b011010111010;
        mem[6817] = 12'b011010111010;
        mem[6818] = 12'b011010111001;
        mem[6819] = 12'b011010111001;
        mem[6820] = 12'b011010111001;
        mem[6821] = 12'b011010111000;
        mem[6822] = 12'b011010111000;
        mem[6823] = 12'b011010111000;
        mem[6824] = 12'b011010110111;
        mem[6825] = 12'b011010110111;
        mem[6826] = 12'b011010110111;
        mem[6827] = 12'b011010110110;
        mem[6828] = 12'b011010110110;
        mem[6829] = 12'b011010110110;
        mem[6830] = 12'b011010110101;
        mem[6831] = 12'b011010110101;
        mem[6832] = 12'b011010110100;
        mem[6833] = 12'b011010110100;
        mem[6834] = 12'b011010110100;
        mem[6835] = 12'b011010110011;
        mem[6836] = 12'b011010110011;
        mem[6837] = 12'b011010110011;
        mem[6838] = 12'b011010110010;
        mem[6839] = 12'b011010110010;
        mem[6840] = 12'b011010110010;
        mem[6841] = 12'b011010110001;
        mem[6842] = 12'b011010110001;
        mem[6843] = 12'b011010110001;
        mem[6844] = 12'b011010110000;
        mem[6845] = 12'b011010110000;
        mem[6846] = 12'b011010110000;
        mem[6847] = 12'b011010101111;
        mem[6848] = 12'b011010101111;
        mem[6849] = 12'b011010101111;
        mem[6850] = 12'b011010101110;
        mem[6851] = 12'b011010101110;
        mem[6852] = 12'b011010101101;
        mem[6853] = 12'b011010101101;
        mem[6854] = 12'b011010101101;
        mem[6855] = 12'b011010101100;
        mem[6856] = 12'b011010101100;
        mem[6857] = 12'b011010101100;
        mem[6858] = 12'b011010101011;
        mem[6859] = 12'b011010101011;
        mem[6860] = 12'b011010101011;
        mem[6861] = 12'b011010101010;
        mem[6862] = 12'b011010101010;
        mem[6863] = 12'b011010101010;
        mem[6864] = 12'b011010101001;
        mem[6865] = 12'b011010101001;
        mem[6866] = 12'b011010101000;
        mem[6867] = 12'b011010101000;
        mem[6868] = 12'b011010101000;
        mem[6869] = 12'b011010100111;
        mem[6870] = 12'b011010100111;
        mem[6871] = 12'b011010100111;
        mem[6872] = 12'b011010100110;
        mem[6873] = 12'b011010100110;
        mem[6874] = 12'b011010100110;
        mem[6875] = 12'b011010100101;
        mem[6876] = 12'b011010100101;
        mem[6877] = 12'b011010100101;
        mem[6878] = 12'b011010100100;
        mem[6879] = 12'b011010100100;
        mem[6880] = 12'b011010100011;
        mem[6881] = 12'b011010100011;
        mem[6882] = 12'b011010100011;
        mem[6883] = 12'b011010100010;
        mem[6884] = 12'b011010100010;
        mem[6885] = 12'b011010100010;
        mem[6886] = 12'b011010100001;
        mem[6887] = 12'b011010100001;
        mem[6888] = 12'b011010100001;
        mem[6889] = 12'b011010100000;
        mem[6890] = 12'b011010100000;
        mem[6891] = 12'b011010100000;
        mem[6892] = 12'b011010011111;
        mem[6893] = 12'b011010011111;
        mem[6894] = 12'b011010011110;
        mem[6895] = 12'b011010011110;
        mem[6896] = 12'b011010011110;
        mem[6897] = 12'b011010011101;
        mem[6898] = 12'b011010011101;
        mem[6899] = 12'b011010011101;
        mem[6900] = 12'b011010011100;
        mem[6901] = 12'b011010011100;
        mem[6902] = 12'b011010011100;
        mem[6903] = 12'b011010011011;
        mem[6904] = 12'b011010011011;
        mem[6905] = 12'b011010011010;
        mem[6906] = 12'b011010011010;
        mem[6907] = 12'b011010011010;
        mem[6908] = 12'b011010011001;
        mem[6909] = 12'b011010011001;
        mem[6910] = 12'b011010011001;
        mem[6911] = 12'b011010011000;
        mem[6912] = 12'b011010011000;
        mem[6913] = 12'b011010011000;
        mem[6914] = 12'b011010010111;
        mem[6915] = 12'b011010010111;
        mem[6916] = 12'b011010010110;
        mem[6917] = 12'b011010010110;
        mem[6918] = 12'b011010010110;
        mem[6919] = 12'b011010010101;
        mem[6920] = 12'b011010010101;
        mem[6921] = 12'b011010010101;
        mem[6922] = 12'b011010010100;
        mem[6923] = 12'b011010010100;
        mem[6924] = 12'b011010010100;
        mem[6925] = 12'b011010010011;
        mem[6926] = 12'b011010010011;
        mem[6927] = 12'b011010010010;
        mem[6928] = 12'b011010010010;
        mem[6929] = 12'b011010010010;
        mem[6930] = 12'b011010010001;
        mem[6931] = 12'b011010010001;
        mem[6932] = 12'b011010010001;
        mem[6933] = 12'b011010010000;
        mem[6934] = 12'b011010010000;
        mem[6935] = 12'b011010010000;
        mem[6936] = 12'b011010001111;
        mem[6937] = 12'b011010001111;
        mem[6938] = 12'b011010001110;
        mem[6939] = 12'b011010001110;
        mem[6940] = 12'b011010001110;
        mem[6941] = 12'b011010001101;
        mem[6942] = 12'b011010001101;
        mem[6943] = 12'b011010001101;
        mem[6944] = 12'b011010001100;
        mem[6945] = 12'b011010001100;
        mem[6946] = 12'b011010001011;
        mem[6947] = 12'b011010001011;
        mem[6948] = 12'b011010001011;
        mem[6949] = 12'b011010001010;
        mem[6950] = 12'b011010001010;
        mem[6951] = 12'b011010001010;
        mem[6952] = 12'b011010001001;
        mem[6953] = 12'b011010001001;
        mem[6954] = 12'b011010001001;
        mem[6955] = 12'b011010001000;
        mem[6956] = 12'b011010001000;
        mem[6957] = 12'b011010000111;
        mem[6958] = 12'b011010000111;
        mem[6959] = 12'b011010000111;
        mem[6960] = 12'b011010000110;
        mem[6961] = 12'b011010000110;
        mem[6962] = 12'b011010000110;
        mem[6963] = 12'b011010000101;
        mem[6964] = 12'b011010000101;
        mem[6965] = 12'b011010000100;
        mem[6966] = 12'b011010000100;
        mem[6967] = 12'b011010000100;
        mem[6968] = 12'b011010000011;
        mem[6969] = 12'b011010000011;
        mem[6970] = 12'b011010000011;
        mem[6971] = 12'b011010000010;
        mem[6972] = 12'b011010000010;
        mem[6973] = 12'b011010000001;
        mem[6974] = 12'b011010000001;
        mem[6975] = 12'b011010000001;
        mem[6976] = 12'b011010000000;
        mem[6977] = 12'b011010000000;
        mem[6978] = 12'b011010000000;
        mem[6979] = 12'b011001111111;
        mem[6980] = 12'b011001111111;
        mem[6981] = 12'b011001111110;
        mem[6982] = 12'b011001111110;
        mem[6983] = 12'b011001111110;
        mem[6984] = 12'b011001111101;
        mem[6985] = 12'b011001111101;
        mem[6986] = 12'b011001111101;
        mem[6987] = 12'b011001111100;
        mem[6988] = 12'b011001111100;
        mem[6989] = 12'b011001111011;
        mem[6990] = 12'b011001111011;
        mem[6991] = 12'b011001111011;
        mem[6992] = 12'b011001111010;
        mem[6993] = 12'b011001111010;
        mem[6994] = 12'b011001111010;
        mem[6995] = 12'b011001111001;
        mem[6996] = 12'b011001111001;
        mem[6997] = 12'b011001111000;
        mem[6998] = 12'b011001111000;
        mem[6999] = 12'b011001111000;
        mem[7000] = 12'b011001110111;
        mem[7001] = 12'b011001110111;
        mem[7002] = 12'b011001110111;
        mem[7003] = 12'b011001110110;
        mem[7004] = 12'b011001110110;
        mem[7005] = 12'b011001110101;
        mem[7006] = 12'b011001110101;
        mem[7007] = 12'b011001110101;
        mem[7008] = 12'b011001110100;
        mem[7009] = 12'b011001110100;
        mem[7010] = 12'b011001110100;
        mem[7011] = 12'b011001110011;
        mem[7012] = 12'b011001110011;
        mem[7013] = 12'b011001110010;
        mem[7014] = 12'b011001110010;
        mem[7015] = 12'b011001110010;
        mem[7016] = 12'b011001110001;
        mem[7017] = 12'b011001110001;
        mem[7018] = 12'b011001110000;
        mem[7019] = 12'b011001110000;
        mem[7020] = 12'b011001110000;
        mem[7021] = 12'b011001101111;
        mem[7022] = 12'b011001101111;
        mem[7023] = 12'b011001101111;
        mem[7024] = 12'b011001101110;
        mem[7025] = 12'b011001101110;
        mem[7026] = 12'b011001101101;
        mem[7027] = 12'b011001101101;
        mem[7028] = 12'b011001101101;
        mem[7029] = 12'b011001101100;
        mem[7030] = 12'b011001101100;
        mem[7031] = 12'b011001101011;
        mem[7032] = 12'b011001101011;
        mem[7033] = 12'b011001101011;
        mem[7034] = 12'b011001101010;
        mem[7035] = 12'b011001101010;
        mem[7036] = 12'b011001101010;
        mem[7037] = 12'b011001101001;
        mem[7038] = 12'b011001101001;
        mem[7039] = 12'b011001101000;
        mem[7040] = 12'b011001101000;
        mem[7041] = 12'b011001101000;
        mem[7042] = 12'b011001100111;
        mem[7043] = 12'b011001100111;
        mem[7044] = 12'b011001100110;
        mem[7045] = 12'b011001100110;
        mem[7046] = 12'b011001100110;
        mem[7047] = 12'b011001100101;
        mem[7048] = 12'b011001100101;
        mem[7049] = 12'b011001100101;
        mem[7050] = 12'b011001100100;
        mem[7051] = 12'b011001100100;
        mem[7052] = 12'b011001100011;
        mem[7053] = 12'b011001100011;
        mem[7054] = 12'b011001100011;
        mem[7055] = 12'b011001100010;
        mem[7056] = 12'b011001100010;
        mem[7057] = 12'b011001100001;
        mem[7058] = 12'b011001100001;
        mem[7059] = 12'b011001100001;
        mem[7060] = 12'b011001100000;
        mem[7061] = 12'b011001100000;
        mem[7062] = 12'b011001100000;
        mem[7063] = 12'b011001011111;
        mem[7064] = 12'b011001011111;
        mem[7065] = 12'b011001011110;
        mem[7066] = 12'b011001011110;
        mem[7067] = 12'b011001011110;
        mem[7068] = 12'b011001011101;
        mem[7069] = 12'b011001011101;
        mem[7070] = 12'b011001011100;
        mem[7071] = 12'b011001011100;
        mem[7072] = 12'b011001011100;
        mem[7073] = 12'b011001011011;
        mem[7074] = 12'b011001011011;
        mem[7075] = 12'b011001011010;
        mem[7076] = 12'b011001011010;
        mem[7077] = 12'b011001011010;
        mem[7078] = 12'b011001011001;
        mem[7079] = 12'b011001011001;
        mem[7080] = 12'b011001011001;
        mem[7081] = 12'b011001011000;
        mem[7082] = 12'b011001011000;
        mem[7083] = 12'b011001010111;
        mem[7084] = 12'b011001010111;
        mem[7085] = 12'b011001010111;
        mem[7086] = 12'b011001010110;
        mem[7087] = 12'b011001010110;
        mem[7088] = 12'b011001010101;
        mem[7089] = 12'b011001010101;
        mem[7090] = 12'b011001010101;
        mem[7091] = 12'b011001010100;
        mem[7092] = 12'b011001010100;
        mem[7093] = 12'b011001010011;
        mem[7094] = 12'b011001010011;
        mem[7095] = 12'b011001010011;
        mem[7096] = 12'b011001010010;
        mem[7097] = 12'b011001010010;
        mem[7098] = 12'b011001010001;
        mem[7099] = 12'b011001010001;
        mem[7100] = 12'b011001010001;
        mem[7101] = 12'b011001010000;
        mem[7102] = 12'b011001010000;
        mem[7103] = 12'b011001001111;
        mem[7104] = 12'b011001001111;
        mem[7105] = 12'b011001001111;
        mem[7106] = 12'b011001001110;
        mem[7107] = 12'b011001001110;
        mem[7108] = 12'b011001001110;
        mem[7109] = 12'b011001001101;
        mem[7110] = 12'b011001001101;
        mem[7111] = 12'b011001001100;
        mem[7112] = 12'b011001001100;
        mem[7113] = 12'b011001001100;
        mem[7114] = 12'b011001001011;
        mem[7115] = 12'b011001001011;
        mem[7116] = 12'b011001001010;
        mem[7117] = 12'b011001001010;
        mem[7118] = 12'b011001001010;
        mem[7119] = 12'b011001001001;
        mem[7120] = 12'b011001001001;
        mem[7121] = 12'b011001001000;
        mem[7122] = 12'b011001001000;
        mem[7123] = 12'b011001001000;
        mem[7124] = 12'b011001000111;
        mem[7125] = 12'b011001000111;
        mem[7126] = 12'b011001000110;
        mem[7127] = 12'b011001000110;
        mem[7128] = 12'b011001000110;
        mem[7129] = 12'b011001000101;
        mem[7130] = 12'b011001000101;
        mem[7131] = 12'b011001000100;
        mem[7132] = 12'b011001000100;
        mem[7133] = 12'b011001000100;
        mem[7134] = 12'b011001000011;
        mem[7135] = 12'b011001000011;
        mem[7136] = 12'b011001000010;
        mem[7137] = 12'b011001000010;
        mem[7138] = 12'b011001000010;
        mem[7139] = 12'b011001000001;
        mem[7140] = 12'b011001000001;
        mem[7141] = 12'b011001000000;
        mem[7142] = 12'b011001000000;
        mem[7143] = 12'b011001000000;
        mem[7144] = 12'b011000111111;
        mem[7145] = 12'b011000111111;
        mem[7146] = 12'b011000111110;
        mem[7147] = 12'b011000111110;
        mem[7148] = 12'b011000111110;
        mem[7149] = 12'b011000111101;
        mem[7150] = 12'b011000111101;
        mem[7151] = 12'b011000111100;
        mem[7152] = 12'b011000111100;
        mem[7153] = 12'b011000111100;
        mem[7154] = 12'b011000111011;
        mem[7155] = 12'b011000111011;
        mem[7156] = 12'b011000111010;
        mem[7157] = 12'b011000111010;
        mem[7158] = 12'b011000111010;
        mem[7159] = 12'b011000111001;
        mem[7160] = 12'b011000111001;
        mem[7161] = 12'b011000111000;
        mem[7162] = 12'b011000111000;
        mem[7163] = 12'b011000111000;
        mem[7164] = 12'b011000110111;
        mem[7165] = 12'b011000110111;
        mem[7166] = 12'b011000110110;
        mem[7167] = 12'b011000110110;
        mem[7168] = 12'b011000110101;
        mem[7169] = 12'b011000110101;
        mem[7170] = 12'b011000110101;
        mem[7171] = 12'b011000110100;
        mem[7172] = 12'b011000110100;
        mem[7173] = 12'b011000110011;
        mem[7174] = 12'b011000110011;
        mem[7175] = 12'b011000110011;
        mem[7176] = 12'b011000110010;
        mem[7177] = 12'b011000110010;
        mem[7178] = 12'b011000110001;
        mem[7179] = 12'b011000110001;
        mem[7180] = 12'b011000110001;
        mem[7181] = 12'b011000110000;
        mem[7182] = 12'b011000110000;
        mem[7183] = 12'b011000101111;
        mem[7184] = 12'b011000101111;
        mem[7185] = 12'b011000101111;
        mem[7186] = 12'b011000101110;
        mem[7187] = 12'b011000101110;
        mem[7188] = 12'b011000101101;
        mem[7189] = 12'b011000101101;
        mem[7190] = 12'b011000101101;
        mem[7191] = 12'b011000101100;
        mem[7192] = 12'b011000101100;
        mem[7193] = 12'b011000101011;
        mem[7194] = 12'b011000101011;
        mem[7195] = 12'b011000101010;
        mem[7196] = 12'b011000101010;
        mem[7197] = 12'b011000101010;
        mem[7198] = 12'b011000101001;
        mem[7199] = 12'b011000101001;
        mem[7200] = 12'b011000101000;
        mem[7201] = 12'b011000101000;
        mem[7202] = 12'b011000101000;
        mem[7203] = 12'b011000100111;
        mem[7204] = 12'b011000100111;
        mem[7205] = 12'b011000100110;
        mem[7206] = 12'b011000100110;
        mem[7207] = 12'b011000100110;
        mem[7208] = 12'b011000100101;
        mem[7209] = 12'b011000100101;
        mem[7210] = 12'b011000100100;
        mem[7211] = 12'b011000100100;
        mem[7212] = 12'b011000100100;
        mem[7213] = 12'b011000100011;
        mem[7214] = 12'b011000100011;
        mem[7215] = 12'b011000100010;
        mem[7216] = 12'b011000100010;
        mem[7217] = 12'b011000100001;
        mem[7218] = 12'b011000100001;
        mem[7219] = 12'b011000100001;
        mem[7220] = 12'b011000100000;
        mem[7221] = 12'b011000100000;
        mem[7222] = 12'b011000011111;
        mem[7223] = 12'b011000011111;
        mem[7224] = 12'b011000011111;
        mem[7225] = 12'b011000011110;
        mem[7226] = 12'b011000011110;
        mem[7227] = 12'b011000011101;
        mem[7228] = 12'b011000011101;
        mem[7229] = 12'b011000011100;
        mem[7230] = 12'b011000011100;
        mem[7231] = 12'b011000011100;
        mem[7232] = 12'b011000011011;
        mem[7233] = 12'b011000011011;
        mem[7234] = 12'b011000011010;
        mem[7235] = 12'b011000011010;
        mem[7236] = 12'b011000011010;
        mem[7237] = 12'b011000011001;
        mem[7238] = 12'b011000011001;
        mem[7239] = 12'b011000011000;
        mem[7240] = 12'b011000011000;
        mem[7241] = 12'b011000011000;
        mem[7242] = 12'b011000010111;
        mem[7243] = 12'b011000010111;
        mem[7244] = 12'b011000010110;
        mem[7245] = 12'b011000010110;
        mem[7246] = 12'b011000010101;
        mem[7247] = 12'b011000010101;
        mem[7248] = 12'b011000010101;
        mem[7249] = 12'b011000010100;
        mem[7250] = 12'b011000010100;
        mem[7251] = 12'b011000010011;
        mem[7252] = 12'b011000010011;
        mem[7253] = 12'b011000010010;
        mem[7254] = 12'b011000010010;
        mem[7255] = 12'b011000010010;
        mem[7256] = 12'b011000010001;
        mem[7257] = 12'b011000010001;
        mem[7258] = 12'b011000010000;
        mem[7259] = 12'b011000010000;
        mem[7260] = 12'b011000010000;
        mem[7261] = 12'b011000001111;
        mem[7262] = 12'b011000001111;
        mem[7263] = 12'b011000001110;
        mem[7264] = 12'b011000001110;
        mem[7265] = 12'b011000001101;
        mem[7266] = 12'b011000001101;
        mem[7267] = 12'b011000001101;
        mem[7268] = 12'b011000001100;
        mem[7269] = 12'b011000001100;
        mem[7270] = 12'b011000001011;
        mem[7271] = 12'b011000001011;
        mem[7272] = 12'b011000001011;
        mem[7273] = 12'b011000001010;
        mem[7274] = 12'b011000001010;
        mem[7275] = 12'b011000001001;
        mem[7276] = 12'b011000001001;
        mem[7277] = 12'b011000001000;
        mem[7278] = 12'b011000001000;
        mem[7279] = 12'b011000001000;
        mem[7280] = 12'b011000000111;
        mem[7281] = 12'b011000000111;
        mem[7282] = 12'b011000000110;
        mem[7283] = 12'b011000000110;
        mem[7284] = 12'b011000000101;
        mem[7285] = 12'b011000000101;
        mem[7286] = 12'b011000000101;
        mem[7287] = 12'b011000000100;
        mem[7288] = 12'b011000000100;
        mem[7289] = 12'b011000000011;
        mem[7290] = 12'b011000000011;
        mem[7291] = 12'b011000000010;
        mem[7292] = 12'b011000000010;
        mem[7293] = 12'b011000000010;
        mem[7294] = 12'b011000000001;
        mem[7295] = 12'b011000000001;
        mem[7296] = 12'b011000000000;
        mem[7297] = 12'b011000000000;
        mem[7298] = 12'b011000000000;
        mem[7299] = 12'b010111111111;
        mem[7300] = 12'b010111111111;
        mem[7301] = 12'b010111111110;
        mem[7302] = 12'b010111111110;
        mem[7303] = 12'b010111111101;
        mem[7304] = 12'b010111111101;
        mem[7305] = 12'b010111111101;
        mem[7306] = 12'b010111111100;
        mem[7307] = 12'b010111111100;
        mem[7308] = 12'b010111111011;
        mem[7309] = 12'b010111111011;
        mem[7310] = 12'b010111111010;
        mem[7311] = 12'b010111111010;
        mem[7312] = 12'b010111111010;
        mem[7313] = 12'b010111111001;
        mem[7314] = 12'b010111111001;
        mem[7315] = 12'b010111111000;
        mem[7316] = 12'b010111111000;
        mem[7317] = 12'b010111110111;
        mem[7318] = 12'b010111110111;
        mem[7319] = 12'b010111110111;
        mem[7320] = 12'b010111110110;
        mem[7321] = 12'b010111110110;
        mem[7322] = 12'b010111110101;
        mem[7323] = 12'b010111110101;
        mem[7324] = 12'b010111110100;
        mem[7325] = 12'b010111110100;
        mem[7326] = 12'b010111110100;
        mem[7327] = 12'b010111110011;
        mem[7328] = 12'b010111110011;
        mem[7329] = 12'b010111110010;
        mem[7330] = 12'b010111110010;
        mem[7331] = 12'b010111110001;
        mem[7332] = 12'b010111110001;
        mem[7333] = 12'b010111110001;
        mem[7334] = 12'b010111110000;
        mem[7335] = 12'b010111110000;
        mem[7336] = 12'b010111101111;
        mem[7337] = 12'b010111101111;
        mem[7338] = 12'b010111101110;
        mem[7339] = 12'b010111101110;
        mem[7340] = 12'b010111101110;
        mem[7341] = 12'b010111101101;
        mem[7342] = 12'b010111101101;
        mem[7343] = 12'b010111101100;
        mem[7344] = 12'b010111101100;
        mem[7345] = 12'b010111101011;
        mem[7346] = 12'b010111101011;
        mem[7347] = 12'b010111101011;
        mem[7348] = 12'b010111101010;
        mem[7349] = 12'b010111101010;
        mem[7350] = 12'b010111101001;
        mem[7351] = 12'b010111101001;
        mem[7352] = 12'b010111101000;
        mem[7353] = 12'b010111101000;
        mem[7354] = 12'b010111100111;
        mem[7355] = 12'b010111100111;
        mem[7356] = 12'b010111100111;
        mem[7357] = 12'b010111100110;
        mem[7358] = 12'b010111100110;
        mem[7359] = 12'b010111100101;
        mem[7360] = 12'b010111100101;
        mem[7361] = 12'b010111100100;
        mem[7362] = 12'b010111100100;
        mem[7363] = 12'b010111100100;
        mem[7364] = 12'b010111100011;
        mem[7365] = 12'b010111100011;
        mem[7366] = 12'b010111100010;
        mem[7367] = 12'b010111100010;
        mem[7368] = 12'b010111100001;
        mem[7369] = 12'b010111100001;
        mem[7370] = 12'b010111100001;
        mem[7371] = 12'b010111100000;
        mem[7372] = 12'b010111100000;
        mem[7373] = 12'b010111011111;
        mem[7374] = 12'b010111011111;
        mem[7375] = 12'b010111011110;
        mem[7376] = 12'b010111011110;
        mem[7377] = 12'b010111011101;
        mem[7378] = 12'b010111011101;
        mem[7379] = 12'b010111011101;
        mem[7380] = 12'b010111011100;
        mem[7381] = 12'b010111011100;
        mem[7382] = 12'b010111011011;
        mem[7383] = 12'b010111011011;
        mem[7384] = 12'b010111011010;
        mem[7385] = 12'b010111011010;
        mem[7386] = 12'b010111011010;
        mem[7387] = 12'b010111011001;
        mem[7388] = 12'b010111011001;
        mem[7389] = 12'b010111011000;
        mem[7390] = 12'b010111011000;
        mem[7391] = 12'b010111010111;
        mem[7392] = 12'b010111010111;
        mem[7393] = 12'b010111010110;
        mem[7394] = 12'b010111010110;
        mem[7395] = 12'b010111010110;
        mem[7396] = 12'b010111010101;
        mem[7397] = 12'b010111010101;
        mem[7398] = 12'b010111010100;
        mem[7399] = 12'b010111010100;
        mem[7400] = 12'b010111010011;
        mem[7401] = 12'b010111010011;
        mem[7402] = 12'b010111010010;
        mem[7403] = 12'b010111010010;
        mem[7404] = 12'b010111010010;
        mem[7405] = 12'b010111010001;
        mem[7406] = 12'b010111010001;
        mem[7407] = 12'b010111010000;
        mem[7408] = 12'b010111010000;
        mem[7409] = 12'b010111001111;
        mem[7410] = 12'b010111001111;
        mem[7411] = 12'b010111001111;
        mem[7412] = 12'b010111001110;
        mem[7413] = 12'b010111001110;
        mem[7414] = 12'b010111001101;
        mem[7415] = 12'b010111001101;
        mem[7416] = 12'b010111001100;
        mem[7417] = 12'b010111001100;
        mem[7418] = 12'b010111001011;
        mem[7419] = 12'b010111001011;
        mem[7420] = 12'b010111001011;
        mem[7421] = 12'b010111001010;
        mem[7422] = 12'b010111001010;
        mem[7423] = 12'b010111001001;
        mem[7424] = 12'b010111001001;
        mem[7425] = 12'b010111001000;
        mem[7426] = 12'b010111001000;
        mem[7427] = 12'b010111000111;
        mem[7428] = 12'b010111000111;
        mem[7429] = 12'b010111000111;
        mem[7430] = 12'b010111000110;
        mem[7431] = 12'b010111000110;
        mem[7432] = 12'b010111000101;
        mem[7433] = 12'b010111000101;
        mem[7434] = 12'b010111000100;
        mem[7435] = 12'b010111000100;
        mem[7436] = 12'b010111000011;
        mem[7437] = 12'b010111000011;
        mem[7438] = 12'b010111000011;
        mem[7439] = 12'b010111000010;
        mem[7440] = 12'b010111000010;
        mem[7441] = 12'b010111000001;
        mem[7442] = 12'b010111000001;
        mem[7443] = 12'b010111000000;
        mem[7444] = 12'b010111000000;
        mem[7445] = 12'b010110111111;
        mem[7446] = 12'b010110111111;
        mem[7447] = 12'b010110111111;
        mem[7448] = 12'b010110111110;
        mem[7449] = 12'b010110111110;
        mem[7450] = 12'b010110111101;
        mem[7451] = 12'b010110111101;
        mem[7452] = 12'b010110111100;
        mem[7453] = 12'b010110111100;
        mem[7454] = 12'b010110111011;
        mem[7455] = 12'b010110111011;
        mem[7456] = 12'b010110111010;
        mem[7457] = 12'b010110111010;
        mem[7458] = 12'b010110111010;
        mem[7459] = 12'b010110111001;
        mem[7460] = 12'b010110111001;
        mem[7461] = 12'b010110111000;
        mem[7462] = 12'b010110111000;
        mem[7463] = 12'b010110110111;
        mem[7464] = 12'b010110110111;
        mem[7465] = 12'b010110110110;
        mem[7466] = 12'b010110110110;
        mem[7467] = 12'b010110110110;
        mem[7468] = 12'b010110110101;
        mem[7469] = 12'b010110110101;
        mem[7470] = 12'b010110110100;
        mem[7471] = 12'b010110110100;
        mem[7472] = 12'b010110110011;
        mem[7473] = 12'b010110110011;
        mem[7474] = 12'b010110110010;
        mem[7475] = 12'b010110110010;
        mem[7476] = 12'b010110110001;
        mem[7477] = 12'b010110110001;
        mem[7478] = 12'b010110110001;
        mem[7479] = 12'b010110110000;
        mem[7480] = 12'b010110110000;
        mem[7481] = 12'b010110101111;
        mem[7482] = 12'b010110101111;
        mem[7483] = 12'b010110101110;
        mem[7484] = 12'b010110101110;
        mem[7485] = 12'b010110101101;
        mem[7486] = 12'b010110101101;
        mem[7487] = 12'b010110101101;
        mem[7488] = 12'b010110101100;
        mem[7489] = 12'b010110101100;
        mem[7490] = 12'b010110101011;
        mem[7491] = 12'b010110101011;
        mem[7492] = 12'b010110101010;
        mem[7493] = 12'b010110101010;
        mem[7494] = 12'b010110101001;
        mem[7495] = 12'b010110101001;
        mem[7496] = 12'b010110101000;
        mem[7497] = 12'b010110101000;
        mem[7498] = 12'b010110101000;
        mem[7499] = 12'b010110100111;
        mem[7500] = 12'b010110100111;
        mem[7501] = 12'b010110100110;
        mem[7502] = 12'b010110100110;
        mem[7503] = 12'b010110100101;
        mem[7504] = 12'b010110100101;
        mem[7505] = 12'b010110100100;
        mem[7506] = 12'b010110100100;
        mem[7507] = 12'b010110100011;
        mem[7508] = 12'b010110100011;
        mem[7509] = 12'b010110100011;
        mem[7510] = 12'b010110100010;
        mem[7511] = 12'b010110100010;
        mem[7512] = 12'b010110100001;
        mem[7513] = 12'b010110100001;
        mem[7514] = 12'b010110100000;
        mem[7515] = 12'b010110100000;
        mem[7516] = 12'b010110011111;
        mem[7517] = 12'b010110011111;
        mem[7518] = 12'b010110011110;
        mem[7519] = 12'b010110011110;
        mem[7520] = 12'b010110011101;
        mem[7521] = 12'b010110011101;
        mem[7522] = 12'b010110011101;
        mem[7523] = 12'b010110011100;
        mem[7524] = 12'b010110011100;
        mem[7525] = 12'b010110011011;
        mem[7526] = 12'b010110011011;
        mem[7527] = 12'b010110011010;
        mem[7528] = 12'b010110011010;
        mem[7529] = 12'b010110011001;
        mem[7530] = 12'b010110011001;
        mem[7531] = 12'b010110011000;
        mem[7532] = 12'b010110011000;
        mem[7533] = 12'b010110011000;
        mem[7534] = 12'b010110010111;
        mem[7535] = 12'b010110010111;
        mem[7536] = 12'b010110010110;
        mem[7537] = 12'b010110010110;
        mem[7538] = 12'b010110010101;
        mem[7539] = 12'b010110010101;
        mem[7540] = 12'b010110010100;
        mem[7541] = 12'b010110010100;
        mem[7542] = 12'b010110010011;
        mem[7543] = 12'b010110010011;
        mem[7544] = 12'b010110010010;
        mem[7545] = 12'b010110010010;
        mem[7546] = 12'b010110010010;
        mem[7547] = 12'b010110010001;
        mem[7548] = 12'b010110010001;
        mem[7549] = 12'b010110010000;
        mem[7550] = 12'b010110010000;
        mem[7551] = 12'b010110001111;
        mem[7552] = 12'b010110001111;
        mem[7553] = 12'b010110001110;
        mem[7554] = 12'b010110001110;
        mem[7555] = 12'b010110001101;
        mem[7556] = 12'b010110001101;
        mem[7557] = 12'b010110001100;
        mem[7558] = 12'b010110001100;
        mem[7559] = 12'b010110001100;
        mem[7560] = 12'b010110001011;
        mem[7561] = 12'b010110001011;
        mem[7562] = 12'b010110001010;
        mem[7563] = 12'b010110001010;
        mem[7564] = 12'b010110001001;
        mem[7565] = 12'b010110001001;
        mem[7566] = 12'b010110001000;
        mem[7567] = 12'b010110001000;
        mem[7568] = 12'b010110000111;
        mem[7569] = 12'b010110000111;
        mem[7570] = 12'b010110000110;
        mem[7571] = 12'b010110000110;
        mem[7572] = 12'b010110000101;
        mem[7573] = 12'b010110000101;
        mem[7574] = 12'b010110000101;
        mem[7575] = 12'b010110000100;
        mem[7576] = 12'b010110000100;
        mem[7577] = 12'b010110000011;
        mem[7578] = 12'b010110000011;
        mem[7579] = 12'b010110000010;
        mem[7580] = 12'b010110000010;
        mem[7581] = 12'b010110000001;
        mem[7582] = 12'b010110000001;
        mem[7583] = 12'b010110000000;
        mem[7584] = 12'b010110000000;
        mem[7585] = 12'b010101111111;
        mem[7586] = 12'b010101111111;
        mem[7587] = 12'b010101111110;
        mem[7588] = 12'b010101111110;
        mem[7589] = 12'b010101111110;
        mem[7590] = 12'b010101111101;
        mem[7591] = 12'b010101111101;
        mem[7592] = 12'b010101111100;
        mem[7593] = 12'b010101111100;
        mem[7594] = 12'b010101111011;
        mem[7595] = 12'b010101111011;
        mem[7596] = 12'b010101111010;
        mem[7597] = 12'b010101111010;
        mem[7598] = 12'b010101111001;
        mem[7599] = 12'b010101111001;
        mem[7600] = 12'b010101111000;
        mem[7601] = 12'b010101111000;
        mem[7602] = 12'b010101110111;
        mem[7603] = 12'b010101110111;
        mem[7604] = 12'b010101110111;
        mem[7605] = 12'b010101110110;
        mem[7606] = 12'b010101110110;
        mem[7607] = 12'b010101110101;
        mem[7608] = 12'b010101110101;
        mem[7609] = 12'b010101110100;
        mem[7610] = 12'b010101110100;
        mem[7611] = 12'b010101110011;
        mem[7612] = 12'b010101110011;
        mem[7613] = 12'b010101110010;
        mem[7614] = 12'b010101110010;
        mem[7615] = 12'b010101110001;
        mem[7616] = 12'b010101110001;
        mem[7617] = 12'b010101110000;
        mem[7618] = 12'b010101110000;
        mem[7619] = 12'b010101101111;
        mem[7620] = 12'b010101101111;
        mem[7621] = 12'b010101101111;
        mem[7622] = 12'b010101101110;
        mem[7623] = 12'b010101101110;
        mem[7624] = 12'b010101101101;
        mem[7625] = 12'b010101101101;
        mem[7626] = 12'b010101101100;
        mem[7627] = 12'b010101101100;
        mem[7628] = 12'b010101101011;
        mem[7629] = 12'b010101101011;
        mem[7630] = 12'b010101101010;
        mem[7631] = 12'b010101101010;
        mem[7632] = 12'b010101101001;
        mem[7633] = 12'b010101101001;
        mem[7634] = 12'b010101101000;
        mem[7635] = 12'b010101101000;
        mem[7636] = 12'b010101100111;
        mem[7637] = 12'b010101100111;
        mem[7638] = 12'b010101100110;
        mem[7639] = 12'b010101100110;
        mem[7640] = 12'b010101100110;
        mem[7641] = 12'b010101100101;
        mem[7642] = 12'b010101100101;
        mem[7643] = 12'b010101100100;
        mem[7644] = 12'b010101100100;
        mem[7645] = 12'b010101100011;
        mem[7646] = 12'b010101100011;
        mem[7647] = 12'b010101100010;
        mem[7648] = 12'b010101100010;
        mem[7649] = 12'b010101100001;
        mem[7650] = 12'b010101100001;
        mem[7651] = 12'b010101100000;
        mem[7652] = 12'b010101100000;
        mem[7653] = 12'b010101011111;
        mem[7654] = 12'b010101011111;
        mem[7655] = 12'b010101011110;
        mem[7656] = 12'b010101011110;
        mem[7657] = 12'b010101011101;
        mem[7658] = 12'b010101011101;
        mem[7659] = 12'b010101011101;
        mem[7660] = 12'b010101011100;
        mem[7661] = 12'b010101011100;
        mem[7662] = 12'b010101011011;
        mem[7663] = 12'b010101011011;
        mem[7664] = 12'b010101011010;
        mem[7665] = 12'b010101011010;
        mem[7666] = 12'b010101011001;
        mem[7667] = 12'b010101011001;
        mem[7668] = 12'b010101011000;
        mem[7669] = 12'b010101011000;
        mem[7670] = 12'b010101010111;
        mem[7671] = 12'b010101010111;
        mem[7672] = 12'b010101010110;
        mem[7673] = 12'b010101010110;
        mem[7674] = 12'b010101010101;
        mem[7675] = 12'b010101010101;
        mem[7676] = 12'b010101010100;
        mem[7677] = 12'b010101010100;
        mem[7678] = 12'b010101010011;
        mem[7679] = 12'b010101010011;
        mem[7680] = 12'b010101010010;
        mem[7681] = 12'b010101010010;
        mem[7682] = 12'b010101010001;
        mem[7683] = 12'b010101010001;
        mem[7684] = 12'b010101010001;
        mem[7685] = 12'b010101010000;
        mem[7686] = 12'b010101010000;
        mem[7687] = 12'b010101001111;
        mem[7688] = 12'b010101001111;
        mem[7689] = 12'b010101001110;
        mem[7690] = 12'b010101001110;
        mem[7691] = 12'b010101001101;
        mem[7692] = 12'b010101001101;
        mem[7693] = 12'b010101001100;
        mem[7694] = 12'b010101001100;
        mem[7695] = 12'b010101001011;
        mem[7696] = 12'b010101001011;
        mem[7697] = 12'b010101001010;
        mem[7698] = 12'b010101001010;
        mem[7699] = 12'b010101001001;
        mem[7700] = 12'b010101001001;
        mem[7701] = 12'b010101001000;
        mem[7702] = 12'b010101001000;
        mem[7703] = 12'b010101000111;
        mem[7704] = 12'b010101000111;
        mem[7705] = 12'b010101000110;
        mem[7706] = 12'b010101000110;
        mem[7707] = 12'b010101000101;
        mem[7708] = 12'b010101000101;
        mem[7709] = 12'b010101000100;
        mem[7710] = 12'b010101000100;
        mem[7711] = 12'b010101000100;
        mem[7712] = 12'b010101000011;
        mem[7713] = 12'b010101000011;
        mem[7714] = 12'b010101000010;
        mem[7715] = 12'b010101000010;
        mem[7716] = 12'b010101000001;
        mem[7717] = 12'b010101000001;
        mem[7718] = 12'b010101000000;
        mem[7719] = 12'b010101000000;
        mem[7720] = 12'b010100111111;
        mem[7721] = 12'b010100111111;
        mem[7722] = 12'b010100111110;
        mem[7723] = 12'b010100111110;
        mem[7724] = 12'b010100111101;
        mem[7725] = 12'b010100111101;
        mem[7726] = 12'b010100111100;
        mem[7727] = 12'b010100111100;
        mem[7728] = 12'b010100111011;
        mem[7729] = 12'b010100111011;
        mem[7730] = 12'b010100111010;
        mem[7731] = 12'b010100111010;
        mem[7732] = 12'b010100111001;
        mem[7733] = 12'b010100111001;
        mem[7734] = 12'b010100111000;
        mem[7735] = 12'b010100111000;
        mem[7736] = 12'b010100110111;
        mem[7737] = 12'b010100110111;
        mem[7738] = 12'b010100110110;
        mem[7739] = 12'b010100110110;
        mem[7740] = 12'b010100110101;
        mem[7741] = 12'b010100110101;
        mem[7742] = 12'b010100110100;
        mem[7743] = 12'b010100110100;
        mem[7744] = 12'b010100110011;
        mem[7745] = 12'b010100110011;
        mem[7746] = 12'b010100110010;
        mem[7747] = 12'b010100110010;
        mem[7748] = 12'b010100110010;
        mem[7749] = 12'b010100110001;
        mem[7750] = 12'b010100110001;
        mem[7751] = 12'b010100110000;
        mem[7752] = 12'b010100110000;
        mem[7753] = 12'b010100101111;
        mem[7754] = 12'b010100101111;
        mem[7755] = 12'b010100101110;
        mem[7756] = 12'b010100101110;
        mem[7757] = 12'b010100101101;
        mem[7758] = 12'b010100101101;
        mem[7759] = 12'b010100101100;
        mem[7760] = 12'b010100101100;
        mem[7761] = 12'b010100101011;
        mem[7762] = 12'b010100101011;
        mem[7763] = 12'b010100101010;
        mem[7764] = 12'b010100101010;
        mem[7765] = 12'b010100101001;
        mem[7766] = 12'b010100101001;
        mem[7767] = 12'b010100101000;
        mem[7768] = 12'b010100101000;
        mem[7769] = 12'b010100100111;
        mem[7770] = 12'b010100100111;
        mem[7771] = 12'b010100100110;
        mem[7772] = 12'b010100100110;
        mem[7773] = 12'b010100100101;
        mem[7774] = 12'b010100100101;
        mem[7775] = 12'b010100100100;
        mem[7776] = 12'b010100100100;
        mem[7777] = 12'b010100100011;
        mem[7778] = 12'b010100100011;
        mem[7779] = 12'b010100100010;
        mem[7780] = 12'b010100100010;
        mem[7781] = 12'b010100100001;
        mem[7782] = 12'b010100100001;
        mem[7783] = 12'b010100100000;
        mem[7784] = 12'b010100100000;
        mem[7785] = 12'b010100011111;
        mem[7786] = 12'b010100011111;
        mem[7787] = 12'b010100011110;
        mem[7788] = 12'b010100011110;
        mem[7789] = 12'b010100011101;
        mem[7790] = 12'b010100011101;
        mem[7791] = 12'b010100011100;
        mem[7792] = 12'b010100011100;
        mem[7793] = 12'b010100011011;
        mem[7794] = 12'b010100011011;
        mem[7795] = 12'b010100011010;
        mem[7796] = 12'b010100011010;
        mem[7797] = 12'b010100011001;
        mem[7798] = 12'b010100011001;
        mem[7799] = 12'b010100011000;
        mem[7800] = 12'b010100011000;
        mem[7801] = 12'b010100010111;
        mem[7802] = 12'b010100010111;
        mem[7803] = 12'b010100010110;
        mem[7804] = 12'b010100010110;
        mem[7805] = 12'b010100010101;
        mem[7806] = 12'b010100010101;
        mem[7807] = 12'b010100010100;
        mem[7808] = 12'b010100010100;
        mem[7809] = 12'b010100010011;
        mem[7810] = 12'b010100010011;
        mem[7811] = 12'b010100010010;
        mem[7812] = 12'b010100010010;
        mem[7813] = 12'b010100010001;
        mem[7814] = 12'b010100010001;
        mem[7815] = 12'b010100010000;
        mem[7816] = 12'b010100010000;
        mem[7817] = 12'b010100001111;
        mem[7818] = 12'b010100001111;
        mem[7819] = 12'b010100001110;
        mem[7820] = 12'b010100001110;
        mem[7821] = 12'b010100001101;
        mem[7822] = 12'b010100001101;
        mem[7823] = 12'b010100001100;
        mem[7824] = 12'b010100001100;
        mem[7825] = 12'b010100001011;
        mem[7826] = 12'b010100001011;
        mem[7827] = 12'b010100001010;
        mem[7828] = 12'b010100001010;
        mem[7829] = 12'b010100001001;
        mem[7830] = 12'b010100001001;
        mem[7831] = 12'b010100001000;
        mem[7832] = 12'b010100001000;
        mem[7833] = 12'b010100000111;
        mem[7834] = 12'b010100000111;
        mem[7835] = 12'b010100000110;
        mem[7836] = 12'b010100000110;
        mem[7837] = 12'b010100000101;
        mem[7838] = 12'b010100000101;
        mem[7839] = 12'b010100000100;
        mem[7840] = 12'b010100000100;
        mem[7841] = 12'b010100000011;
        mem[7842] = 12'b010100000011;
        mem[7843] = 12'b010100000010;
        mem[7844] = 12'b010100000010;
        mem[7845] = 12'b010100000001;
        mem[7846] = 12'b010100000001;
        mem[7847] = 12'b010100000000;
        mem[7848] = 12'b010100000000;
        mem[7849] = 12'b010011111111;
        mem[7850] = 12'b010011111111;
        mem[7851] = 12'b010011111110;
        mem[7852] = 12'b010011111110;
        mem[7853] = 12'b010011111101;
        mem[7854] = 12'b010011111101;
        mem[7855] = 12'b010011111100;
        mem[7856] = 12'b010011111100;
        mem[7857] = 12'b010011111011;
        mem[7858] = 12'b010011111011;
        mem[7859] = 12'b010011111010;
        mem[7860] = 12'b010011111010;
        mem[7861] = 12'b010011111001;
        mem[7862] = 12'b010011111001;
        mem[7863] = 12'b010011111000;
        mem[7864] = 12'b010011111000;
        mem[7865] = 12'b010011110111;
        mem[7866] = 12'b010011110111;
        mem[7867] = 12'b010011110110;
        mem[7868] = 12'b010011110110;
        mem[7869] = 12'b010011110101;
        mem[7870] = 12'b010011110101;
        mem[7871] = 12'b010011110100;
        mem[7872] = 12'b010011110100;
        mem[7873] = 12'b010011110011;
        mem[7874] = 12'b010011110011;
        mem[7875] = 12'b010011110010;
        mem[7876] = 12'b010011110010;
        mem[7877] = 12'b010011110001;
        mem[7878] = 12'b010011110001;
        mem[7879] = 12'b010011110000;
        mem[7880] = 12'b010011110000;
        mem[7881] = 12'b010011101111;
        mem[7882] = 12'b010011101111;
        mem[7883] = 12'b010011101110;
        mem[7884] = 12'b010011101110;
        mem[7885] = 12'b010011101101;
        mem[7886] = 12'b010011101101;
        mem[7887] = 12'b010011101100;
        mem[7888] = 12'b010011101100;
        mem[7889] = 12'b010011101011;
        mem[7890] = 12'b010011101011;
        mem[7891] = 12'b010011101010;
        mem[7892] = 12'b010011101010;
        mem[7893] = 12'b010011101001;
        mem[7894] = 12'b010011101001;
        mem[7895] = 12'b010011101000;
        mem[7896] = 12'b010011101000;
        mem[7897] = 12'b010011100111;
        mem[7898] = 12'b010011100111;
        mem[7899] = 12'b010011100110;
        mem[7900] = 12'b010011100110;
        mem[7901] = 12'b010011100101;
        mem[7902] = 12'b010011100101;
        mem[7903] = 12'b010011100100;
        mem[7904] = 12'b010011100100;
        mem[7905] = 12'b010011100011;
        mem[7906] = 12'b010011100011;
        mem[7907] = 12'b010011100010;
        mem[7908] = 12'b010011100010;
        mem[7909] = 12'b010011100001;
        mem[7910] = 12'b010011100001;
        mem[7911] = 12'b010011100000;
        mem[7912] = 12'b010011100000;
        mem[7913] = 12'b010011011111;
        mem[7914] = 12'b010011011111;
        mem[7915] = 12'b010011011110;
        mem[7916] = 12'b010011011110;
        mem[7917] = 12'b010011011101;
        mem[7918] = 12'b010011011101;
        mem[7919] = 12'b010011011100;
        mem[7920] = 12'b010011011100;
        mem[7921] = 12'b010011011011;
        mem[7922] = 12'b010011011011;
        mem[7923] = 12'b010011011010;
        mem[7924] = 12'b010011011001;
        mem[7925] = 12'b010011011001;
        mem[7926] = 12'b010011011000;
        mem[7927] = 12'b010011011000;
        mem[7928] = 12'b010011010111;
        mem[7929] = 12'b010011010111;
        mem[7930] = 12'b010011010110;
        mem[7931] = 12'b010011010110;
        mem[7932] = 12'b010011010101;
        mem[7933] = 12'b010011010101;
        mem[7934] = 12'b010011010100;
        mem[7935] = 12'b010011010100;
        mem[7936] = 12'b010011010011;
        mem[7937] = 12'b010011010011;
        mem[7938] = 12'b010011010010;
        mem[7939] = 12'b010011010010;
        mem[7940] = 12'b010011010001;
        mem[7941] = 12'b010011010001;
        mem[7942] = 12'b010011010000;
        mem[7943] = 12'b010011010000;
        mem[7944] = 12'b010011001111;
        mem[7945] = 12'b010011001111;
        mem[7946] = 12'b010011001110;
        mem[7947] = 12'b010011001110;
        mem[7948] = 12'b010011001101;
        mem[7949] = 12'b010011001101;
        mem[7950] = 12'b010011001100;
        mem[7951] = 12'b010011001100;
        mem[7952] = 12'b010011001011;
        mem[7953] = 12'b010011001011;
        mem[7954] = 12'b010011001010;
        mem[7955] = 12'b010011001010;
        mem[7956] = 12'b010011001001;
        mem[7957] = 12'b010011001001;
        mem[7958] = 12'b010011001000;
        mem[7959] = 12'b010011001000;
        mem[7960] = 12'b010011000111;
        mem[7961] = 12'b010011000110;
        mem[7962] = 12'b010011000110;
        mem[7963] = 12'b010011000101;
        mem[7964] = 12'b010011000101;
        mem[7965] = 12'b010011000100;
        mem[7966] = 12'b010011000100;
        mem[7967] = 12'b010011000011;
        mem[7968] = 12'b010011000011;
        mem[7969] = 12'b010011000010;
        mem[7970] = 12'b010011000010;
        mem[7971] = 12'b010011000001;
        mem[7972] = 12'b010011000001;
        mem[7973] = 12'b010011000000;
        mem[7974] = 12'b010011000000;
        mem[7975] = 12'b010010111111;
        mem[7976] = 12'b010010111111;
        mem[7977] = 12'b010010111110;
        mem[7978] = 12'b010010111110;
        mem[7979] = 12'b010010111101;
        mem[7980] = 12'b010010111101;
        mem[7981] = 12'b010010111100;
        mem[7982] = 12'b010010111100;
        mem[7983] = 12'b010010111011;
        mem[7984] = 12'b010010111011;
        mem[7985] = 12'b010010111010;
        mem[7986] = 12'b010010111010;
        mem[7987] = 12'b010010111001;
        mem[7988] = 12'b010010111001;
        mem[7989] = 12'b010010111000;
        mem[7990] = 12'b010010110111;
        mem[7991] = 12'b010010110111;
        mem[7992] = 12'b010010110110;
        mem[7993] = 12'b010010110110;
        mem[7994] = 12'b010010110101;
        mem[7995] = 12'b010010110101;
        mem[7996] = 12'b010010110100;
        mem[7997] = 12'b010010110100;
        mem[7998] = 12'b010010110011;
        mem[7999] = 12'b010010110011;
        mem[8000] = 12'b010010110010;
        mem[8001] = 12'b010010110010;
        mem[8002] = 12'b010010110001;
        mem[8003] = 12'b010010110001;
        mem[8004] = 12'b010010110000;
        mem[8005] = 12'b010010110000;
        mem[8006] = 12'b010010101111;
        mem[8007] = 12'b010010101111;
        mem[8008] = 12'b010010101110;
        mem[8009] = 12'b010010101110;
        mem[8010] = 12'b010010101101;
        mem[8011] = 12'b010010101101;
        mem[8012] = 12'b010010101100;
        mem[8013] = 12'b010010101100;
        mem[8014] = 12'b010010101011;
        mem[8015] = 12'b010010101010;
        mem[8016] = 12'b010010101010;
        mem[8017] = 12'b010010101001;
        mem[8018] = 12'b010010101001;
        mem[8019] = 12'b010010101000;
        mem[8020] = 12'b010010101000;
        mem[8021] = 12'b010010100111;
        mem[8022] = 12'b010010100111;
        mem[8023] = 12'b010010100110;
        mem[8024] = 12'b010010100110;
        mem[8025] = 12'b010010100101;
        mem[8026] = 12'b010010100101;
        mem[8027] = 12'b010010100100;
        mem[8028] = 12'b010010100100;
        mem[8029] = 12'b010010100011;
        mem[8030] = 12'b010010100011;
        mem[8031] = 12'b010010100010;
        mem[8032] = 12'b010010100010;
        mem[8033] = 12'b010010100001;
        mem[8034] = 12'b010010100001;
        mem[8035] = 12'b010010100000;
        mem[8036] = 12'b010010011111;
        mem[8037] = 12'b010010011111;
        mem[8038] = 12'b010010011110;
        mem[8039] = 12'b010010011110;
        mem[8040] = 12'b010010011101;
        mem[8041] = 12'b010010011101;
        mem[8042] = 12'b010010011100;
        mem[8043] = 12'b010010011100;
        mem[8044] = 12'b010010011011;
        mem[8045] = 12'b010010011011;
        mem[8046] = 12'b010010011010;
        mem[8047] = 12'b010010011010;
        mem[8048] = 12'b010010011001;
        mem[8049] = 12'b010010011001;
        mem[8050] = 12'b010010011000;
        mem[8051] = 12'b010010011000;
        mem[8052] = 12'b010010010111;
        mem[8053] = 12'b010010010111;
        mem[8054] = 12'b010010010110;
        mem[8055] = 12'b010010010101;
        mem[8056] = 12'b010010010101;
        mem[8057] = 12'b010010010100;
        mem[8058] = 12'b010010010100;
        mem[8059] = 12'b010010010011;
        mem[8060] = 12'b010010010011;
        mem[8061] = 12'b010010010010;
        mem[8062] = 12'b010010010010;
        mem[8063] = 12'b010010010001;
        mem[8064] = 12'b010010010001;
        mem[8065] = 12'b010010010000;
        mem[8066] = 12'b010010010000;
        mem[8067] = 12'b010010001111;
        mem[8068] = 12'b010010001111;
        mem[8069] = 12'b010010001110;
        mem[8070] = 12'b010010001110;
        mem[8071] = 12'b010010001101;
        mem[8072] = 12'b010010001101;
        mem[8073] = 12'b010010001100;
        mem[8074] = 12'b010010001011;
        mem[8075] = 12'b010010001011;
        mem[8076] = 12'b010010001010;
        mem[8077] = 12'b010010001010;
        mem[8078] = 12'b010010001001;
        mem[8079] = 12'b010010001001;
        mem[8080] = 12'b010010001000;
        mem[8081] = 12'b010010001000;
        mem[8082] = 12'b010010000111;
        mem[8083] = 12'b010010000111;
        mem[8084] = 12'b010010000110;
        mem[8085] = 12'b010010000110;
        mem[8086] = 12'b010010000101;
        mem[8087] = 12'b010010000101;
        mem[8088] = 12'b010010000100;
        mem[8089] = 12'b010010000011;
        mem[8090] = 12'b010010000011;
        mem[8091] = 12'b010010000010;
        mem[8092] = 12'b010010000010;
        mem[8093] = 12'b010010000001;
        mem[8094] = 12'b010010000001;
        mem[8095] = 12'b010010000000;
        mem[8096] = 12'b010010000000;
        mem[8097] = 12'b010001111111;
        mem[8098] = 12'b010001111111;
        mem[8099] = 12'b010001111110;
        mem[8100] = 12'b010001111110;
        mem[8101] = 12'b010001111101;
        mem[8102] = 12'b010001111101;
        mem[8103] = 12'b010001111100;
        mem[8104] = 12'b010001111100;
        mem[8105] = 12'b010001111011;
        mem[8106] = 12'b010001111010;
        mem[8107] = 12'b010001111010;
        mem[8108] = 12'b010001111001;
        mem[8109] = 12'b010001111001;
        mem[8110] = 12'b010001111000;
        mem[8111] = 12'b010001111000;
        mem[8112] = 12'b010001110111;
        mem[8113] = 12'b010001110111;
        mem[8114] = 12'b010001110110;
        mem[8115] = 12'b010001110110;
        mem[8116] = 12'b010001110101;
        mem[8117] = 12'b010001110101;
        mem[8118] = 12'b010001110100;
        mem[8119] = 12'b010001110100;
        mem[8120] = 12'b010001110011;
        mem[8121] = 12'b010001110010;
        mem[8122] = 12'b010001110010;
        mem[8123] = 12'b010001110001;
        mem[8124] = 12'b010001110001;
        mem[8125] = 12'b010001110000;
        mem[8126] = 12'b010001110000;
        mem[8127] = 12'b010001101111;
        mem[8128] = 12'b010001101111;
        mem[8129] = 12'b010001101110;
        mem[8130] = 12'b010001101110;
        mem[8131] = 12'b010001101101;
        mem[8132] = 12'b010001101101;
        mem[8133] = 12'b010001101100;
        mem[8134] = 12'b010001101011;
        mem[8135] = 12'b010001101011;
        mem[8136] = 12'b010001101010;
        mem[8137] = 12'b010001101010;
        mem[8138] = 12'b010001101001;
        mem[8139] = 12'b010001101001;
        mem[8140] = 12'b010001101000;
        mem[8141] = 12'b010001101000;
        mem[8142] = 12'b010001100111;
        mem[8143] = 12'b010001100111;
        mem[8144] = 12'b010001100110;
        mem[8145] = 12'b010001100110;
        mem[8146] = 12'b010001100101;
        mem[8147] = 12'b010001100101;
        mem[8148] = 12'b010001100100;
        mem[8149] = 12'b010001100011;
        mem[8150] = 12'b010001100011;
        mem[8151] = 12'b010001100010;
        mem[8152] = 12'b010001100010;
        mem[8153] = 12'b010001100001;
        mem[8154] = 12'b010001100001;
        mem[8155] = 12'b010001100000;
        mem[8156] = 12'b010001100000;
        mem[8157] = 12'b010001011111;
        mem[8158] = 12'b010001011111;
        mem[8159] = 12'b010001011110;
        mem[8160] = 12'b010001011110;
        mem[8161] = 12'b010001011101;
        mem[8162] = 12'b010001011100;
        mem[8163] = 12'b010001011100;
        mem[8164] = 12'b010001011011;
        mem[8165] = 12'b010001011011;
        mem[8166] = 12'b010001011010;
        mem[8167] = 12'b010001011010;
        mem[8168] = 12'b010001011001;
        mem[8169] = 12'b010001011001;
        mem[8170] = 12'b010001011000;
        mem[8171] = 12'b010001011000;
        mem[8172] = 12'b010001010111;
        mem[8173] = 12'b010001010111;
        mem[8174] = 12'b010001010110;
        mem[8175] = 12'b010001010101;
        mem[8176] = 12'b010001010101;
        mem[8177] = 12'b010001010100;
        mem[8178] = 12'b010001010100;
        mem[8179] = 12'b010001010011;
        mem[8180] = 12'b010001010011;
        mem[8181] = 12'b010001010010;
        mem[8182] = 12'b010001010010;
        mem[8183] = 12'b010001010001;
        mem[8184] = 12'b010001010001;
        mem[8185] = 12'b010001010000;
        mem[8186] = 12'b010001001111;
        mem[8187] = 12'b010001001111;
        mem[8188] = 12'b010001001110;
        mem[8189] = 12'b010001001110;
        mem[8190] = 12'b010001001101;
        mem[8191] = 12'b010001001101;
        mem[8192] = 12'b010001001100;
        mem[8193] = 12'b010001001100;
        mem[8194] = 12'b010001001011;
        mem[8195] = 12'b010001001011;
        mem[8196] = 12'b010001001010;
        mem[8197] = 12'b010001001010;
        mem[8198] = 12'b010001001001;
        mem[8199] = 12'b010001001000;
        mem[8200] = 12'b010001001000;
        mem[8201] = 12'b010001000111;
        mem[8202] = 12'b010001000111;
        mem[8203] = 12'b010001000110;
        mem[8204] = 12'b010001000110;
        mem[8205] = 12'b010001000101;
        mem[8206] = 12'b010001000101;
        mem[8207] = 12'b010001000100;
        mem[8208] = 12'b010001000100;
        mem[8209] = 12'b010001000011;
        mem[8210] = 12'b010001000010;
        mem[8211] = 12'b010001000010;
        mem[8212] = 12'b010001000001;
        mem[8213] = 12'b010001000001;
        mem[8214] = 12'b010001000000;
        mem[8215] = 12'b010001000000;
        mem[8216] = 12'b010000111111;
        mem[8217] = 12'b010000111111;
        mem[8218] = 12'b010000111110;
        mem[8219] = 12'b010000111110;
        mem[8220] = 12'b010000111101;
        mem[8221] = 12'b010000111100;
        mem[8222] = 12'b010000111100;
        mem[8223] = 12'b010000111011;
        mem[8224] = 12'b010000111011;
        mem[8225] = 12'b010000111010;
        mem[8226] = 12'b010000111010;
        mem[8227] = 12'b010000111001;
        mem[8228] = 12'b010000111001;
        mem[8229] = 12'b010000111000;
        mem[8230] = 12'b010000111000;
        mem[8231] = 12'b010000110111;
        mem[8232] = 12'b010000110110;
        mem[8233] = 12'b010000110110;
        mem[8234] = 12'b010000110101;
        mem[8235] = 12'b010000110101;
        mem[8236] = 12'b010000110100;
        mem[8237] = 12'b010000110100;
        mem[8238] = 12'b010000110011;
        mem[8239] = 12'b010000110011;
        mem[8240] = 12'b010000110010;
        mem[8241] = 12'b010000110010;
        mem[8242] = 12'b010000110001;
        mem[8243] = 12'b010000110000;
        mem[8244] = 12'b010000110000;
        mem[8245] = 12'b010000101111;
        mem[8246] = 12'b010000101111;
        mem[8247] = 12'b010000101110;
        mem[8248] = 12'b010000101110;
        mem[8249] = 12'b010000101101;
        mem[8250] = 12'b010000101101;
        mem[8251] = 12'b010000101100;
        mem[8252] = 12'b010000101100;
        mem[8253] = 12'b010000101011;
        mem[8254] = 12'b010000101010;
        mem[8255] = 12'b010000101010;
        mem[8256] = 12'b010000101001;
        mem[8257] = 12'b010000101001;
        mem[8258] = 12'b010000101000;
        mem[8259] = 12'b010000101000;
        mem[8260] = 12'b010000100111;
        mem[8261] = 12'b010000100111;
        mem[8262] = 12'b010000100110;
        mem[8263] = 12'b010000100101;
        mem[8264] = 12'b010000100101;
        mem[8265] = 12'b010000100100;
        mem[8266] = 12'b010000100100;
        mem[8267] = 12'b010000100011;
        mem[8268] = 12'b010000100011;
        mem[8269] = 12'b010000100010;
        mem[8270] = 12'b010000100010;
        mem[8271] = 12'b010000100001;
        mem[8272] = 12'b010000100001;
        mem[8273] = 12'b010000100000;
        mem[8274] = 12'b010000011111;
        mem[8275] = 12'b010000011111;
        mem[8276] = 12'b010000011110;
        mem[8277] = 12'b010000011110;
        mem[8278] = 12'b010000011101;
        mem[8279] = 12'b010000011101;
        mem[8280] = 12'b010000011100;
        mem[8281] = 12'b010000011100;
        mem[8282] = 12'b010000011011;
        mem[8283] = 12'b010000011010;
        mem[8284] = 12'b010000011010;
        mem[8285] = 12'b010000011001;
        mem[8286] = 12'b010000011001;
        mem[8287] = 12'b010000011000;
        mem[8288] = 12'b010000011000;
        mem[8289] = 12'b010000010111;
        mem[8290] = 12'b010000010111;
        mem[8291] = 12'b010000010110;
        mem[8292] = 12'b010000010101;
        mem[8293] = 12'b010000010101;
        mem[8294] = 12'b010000010100;
        mem[8295] = 12'b010000010100;
        mem[8296] = 12'b010000010011;
        mem[8297] = 12'b010000010011;
        mem[8298] = 12'b010000010010;
        mem[8299] = 12'b010000010010;
        mem[8300] = 12'b010000010001;
        mem[8301] = 12'b010000010000;
        mem[8302] = 12'b010000010000;
        mem[8303] = 12'b010000001111;
        mem[8304] = 12'b010000001111;
        mem[8305] = 12'b010000001110;
        mem[8306] = 12'b010000001110;
        mem[8307] = 12'b010000001101;
        mem[8308] = 12'b010000001101;
        mem[8309] = 12'b010000001100;
        mem[8310] = 12'b010000001100;
        mem[8311] = 12'b010000001011;
        mem[8312] = 12'b010000001010;
        mem[8313] = 12'b010000001010;
        mem[8314] = 12'b010000001001;
        mem[8315] = 12'b010000001001;
        mem[8316] = 12'b010000001000;
        mem[8317] = 12'b010000001000;
        mem[8318] = 12'b010000000111;
        mem[8319] = 12'b010000000111;
        mem[8320] = 12'b010000000110;
        mem[8321] = 12'b010000000101;
        mem[8322] = 12'b010000000101;
        mem[8323] = 12'b010000000100;
        mem[8324] = 12'b010000000100;
        mem[8325] = 12'b010000000011;
        mem[8326] = 12'b010000000011;
        mem[8327] = 12'b010000000010;
        mem[8328] = 12'b010000000010;
        mem[8329] = 12'b010000000001;
        mem[8330] = 12'b010000000000;
        mem[8331] = 12'b010000000000;
        mem[8332] = 12'b001111111111;
        mem[8333] = 12'b001111111111;
        mem[8334] = 12'b001111111110;
        mem[8335] = 12'b001111111110;
        mem[8336] = 12'b001111111101;
        mem[8337] = 12'b001111111100;
        mem[8338] = 12'b001111111100;
        mem[8339] = 12'b001111111011;
        mem[8340] = 12'b001111111011;
        mem[8341] = 12'b001111111010;
        mem[8342] = 12'b001111111010;
        mem[8343] = 12'b001111111001;
        mem[8344] = 12'b001111111001;
        mem[8345] = 12'b001111111000;
        mem[8346] = 12'b001111110111;
        mem[8347] = 12'b001111110111;
        mem[8348] = 12'b001111110110;
        mem[8349] = 12'b001111110110;
        mem[8350] = 12'b001111110101;
        mem[8351] = 12'b001111110101;
        mem[8352] = 12'b001111110100;
        mem[8353] = 12'b001111110100;
        mem[8354] = 12'b001111110011;
        mem[8355] = 12'b001111110010;
        mem[8356] = 12'b001111110010;
        mem[8357] = 12'b001111110001;
        mem[8358] = 12'b001111110001;
        mem[8359] = 12'b001111110000;
        mem[8360] = 12'b001111110000;
        mem[8361] = 12'b001111101111;
        mem[8362] = 12'b001111101111;
        mem[8363] = 12'b001111101110;
        mem[8364] = 12'b001111101101;
        mem[8365] = 12'b001111101101;
        mem[8366] = 12'b001111101100;
        mem[8367] = 12'b001111101100;
        mem[8368] = 12'b001111101011;
        mem[8369] = 12'b001111101011;
        mem[8370] = 12'b001111101010;
        mem[8371] = 12'b001111101001;
        mem[8372] = 12'b001111101001;
        mem[8373] = 12'b001111101000;
        mem[8374] = 12'b001111101000;
        mem[8375] = 12'b001111100111;
        mem[8376] = 12'b001111100111;
        mem[8377] = 12'b001111100110;
        mem[8378] = 12'b001111100110;
        mem[8379] = 12'b001111100101;
        mem[8380] = 12'b001111100100;
        mem[8381] = 12'b001111100100;
        mem[8382] = 12'b001111100011;
        mem[8383] = 12'b001111100011;
        mem[8384] = 12'b001111100010;
        mem[8385] = 12'b001111100010;
        mem[8386] = 12'b001111100001;
        mem[8387] = 12'b001111100000;
        mem[8388] = 12'b001111100000;
        mem[8389] = 12'b001111011111;
        mem[8390] = 12'b001111011111;
        mem[8391] = 12'b001111011110;
        mem[8392] = 12'b001111011110;
        mem[8393] = 12'b001111011101;
        mem[8394] = 12'b001111011101;
        mem[8395] = 12'b001111011100;
        mem[8396] = 12'b001111011011;
        mem[8397] = 12'b001111011011;
        mem[8398] = 12'b001111011010;
        mem[8399] = 12'b001111011010;
        mem[8400] = 12'b001111011001;
        mem[8401] = 12'b001111011001;
        mem[8402] = 12'b001111011000;
        mem[8403] = 12'b001111010111;
        mem[8404] = 12'b001111010111;
        mem[8405] = 12'b001111010110;
        mem[8406] = 12'b001111010110;
        mem[8407] = 12'b001111010101;
        mem[8408] = 12'b001111010101;
        mem[8409] = 12'b001111010100;
        mem[8410] = 12'b001111010100;
        mem[8411] = 12'b001111010011;
        mem[8412] = 12'b001111010010;
        mem[8413] = 12'b001111010010;
        mem[8414] = 12'b001111010001;
        mem[8415] = 12'b001111010001;
        mem[8416] = 12'b001111010000;
        mem[8417] = 12'b001111010000;
        mem[8418] = 12'b001111001111;
        mem[8419] = 12'b001111001110;
        mem[8420] = 12'b001111001110;
        mem[8421] = 12'b001111001101;
        mem[8422] = 12'b001111001101;
        mem[8423] = 12'b001111001100;
        mem[8424] = 12'b001111001100;
        mem[8425] = 12'b001111001011;
        mem[8426] = 12'b001111001010;
        mem[8427] = 12'b001111001010;
        mem[8428] = 12'b001111001001;
        mem[8429] = 12'b001111001001;
        mem[8430] = 12'b001111001000;
        mem[8431] = 12'b001111001000;
        mem[8432] = 12'b001111000111;
        mem[8433] = 12'b001111000111;
        mem[8434] = 12'b001111000110;
        mem[8435] = 12'b001111000101;
        mem[8436] = 12'b001111000101;
        mem[8437] = 12'b001111000100;
        mem[8438] = 12'b001111000100;
        mem[8439] = 12'b001111000011;
        mem[8440] = 12'b001111000011;
        mem[8441] = 12'b001111000010;
        mem[8442] = 12'b001111000001;
        mem[8443] = 12'b001111000001;
        mem[8444] = 12'b001111000000;
        mem[8445] = 12'b001111000000;
        mem[8446] = 12'b001110111111;
        mem[8447] = 12'b001110111111;
        mem[8448] = 12'b001110111110;
        mem[8449] = 12'b001110111101;
        mem[8450] = 12'b001110111101;
        mem[8451] = 12'b001110111100;
        mem[8452] = 12'b001110111100;
        mem[8453] = 12'b001110111011;
        mem[8454] = 12'b001110111011;
        mem[8455] = 12'b001110111010;
        mem[8456] = 12'b001110111001;
        mem[8457] = 12'b001110111001;
        mem[8458] = 12'b001110111000;
        mem[8459] = 12'b001110111000;
        mem[8460] = 12'b001110110111;
        mem[8461] = 12'b001110110111;
        mem[8462] = 12'b001110110110;
        mem[8463] = 12'b001110110101;
        mem[8464] = 12'b001110110101;
        mem[8465] = 12'b001110110100;
        mem[8466] = 12'b001110110100;
        mem[8467] = 12'b001110110011;
        mem[8468] = 12'b001110110011;
        mem[8469] = 12'b001110110010;
        mem[8470] = 12'b001110110001;
        mem[8471] = 12'b001110110001;
        mem[8472] = 12'b001110110000;
        mem[8473] = 12'b001110110000;
        mem[8474] = 12'b001110101111;
        mem[8475] = 12'b001110101111;
        mem[8476] = 12'b001110101110;
        mem[8477] = 12'b001110101101;
        mem[8478] = 12'b001110101101;
        mem[8479] = 12'b001110101100;
        mem[8480] = 12'b001110101100;
        mem[8481] = 12'b001110101011;
        mem[8482] = 12'b001110101011;
        mem[8483] = 12'b001110101010;
        mem[8484] = 12'b001110101001;
        mem[8485] = 12'b001110101001;
        mem[8486] = 12'b001110101000;
        mem[8487] = 12'b001110101000;
        mem[8488] = 12'b001110100111;
        mem[8489] = 12'b001110100111;
        mem[8490] = 12'b001110100110;
        mem[8491] = 12'b001110100101;
        mem[8492] = 12'b001110100101;
        mem[8493] = 12'b001110100100;
        mem[8494] = 12'b001110100100;
        mem[8495] = 12'b001110100011;
        mem[8496] = 12'b001110100011;
        mem[8497] = 12'b001110100010;
        mem[8498] = 12'b001110100001;
        mem[8499] = 12'b001110100001;
        mem[8500] = 12'b001110100000;
        mem[8501] = 12'b001110100000;
        mem[8502] = 12'b001110011111;
        mem[8503] = 12'b001110011111;
        mem[8504] = 12'b001110011110;
        mem[8505] = 12'b001110011101;
        mem[8506] = 12'b001110011101;
        mem[8507] = 12'b001110011100;
        mem[8508] = 12'b001110011100;
        mem[8509] = 12'b001110011011;
        mem[8510] = 12'b001110011011;
        mem[8511] = 12'b001110011010;
        mem[8512] = 12'b001110011001;
        mem[8513] = 12'b001110011001;
        mem[8514] = 12'b001110011000;
        mem[8515] = 12'b001110011000;
        mem[8516] = 12'b001110010111;
        mem[8517] = 12'b001110010111;
        mem[8518] = 12'b001110010110;
        mem[8519] = 12'b001110010101;
        mem[8520] = 12'b001110010101;
        mem[8521] = 12'b001110010100;
        mem[8522] = 12'b001110010100;
        mem[8523] = 12'b001110010011;
        mem[8524] = 12'b001110010011;
        mem[8525] = 12'b001110010010;
        mem[8526] = 12'b001110010001;
        mem[8527] = 12'b001110010001;
        mem[8528] = 12'b001110010000;
        mem[8529] = 12'b001110010000;
        mem[8530] = 12'b001110001111;
        mem[8531] = 12'b001110001111;
        mem[8532] = 12'b001110001110;
        mem[8533] = 12'b001110001101;
        mem[8534] = 12'b001110001101;
        mem[8535] = 12'b001110001100;
        mem[8536] = 12'b001110001100;
        mem[8537] = 12'b001110001011;
        mem[8538] = 12'b001110001010;
        mem[8539] = 12'b001110001010;
        mem[8540] = 12'b001110001001;
        mem[8541] = 12'b001110001001;
        mem[8542] = 12'b001110001000;
        mem[8543] = 12'b001110001000;
        mem[8544] = 12'b001110000111;
        mem[8545] = 12'b001110000110;
        mem[8546] = 12'b001110000110;
        mem[8547] = 12'b001110000101;
        mem[8548] = 12'b001110000101;
        mem[8549] = 12'b001110000100;
        mem[8550] = 12'b001110000100;
        mem[8551] = 12'b001110000011;
        mem[8552] = 12'b001110000010;
        mem[8553] = 12'b001110000010;
        mem[8554] = 12'b001110000001;
        mem[8555] = 12'b001110000001;
        mem[8556] = 12'b001110000000;
        mem[8557] = 12'b001110000000;
        mem[8558] = 12'b001101111111;
        mem[8559] = 12'b001101111110;
        mem[8560] = 12'b001101111110;
        mem[8561] = 12'b001101111101;
        mem[8562] = 12'b001101111101;
        mem[8563] = 12'b001101111100;
        mem[8564] = 12'b001101111011;
        mem[8565] = 12'b001101111011;
        mem[8566] = 12'b001101111010;
        mem[8567] = 12'b001101111010;
        mem[8568] = 12'b001101111001;
        mem[8569] = 12'b001101111001;
        mem[8570] = 12'b001101111000;
        mem[8571] = 12'b001101110111;
        mem[8572] = 12'b001101110111;
        mem[8573] = 12'b001101110110;
        mem[8574] = 12'b001101110110;
        mem[8575] = 12'b001101110101;
        mem[8576] = 12'b001101110101;
        mem[8577] = 12'b001101110100;
        mem[8578] = 12'b001101110011;
        mem[8579] = 12'b001101110011;
        mem[8580] = 12'b001101110010;
        mem[8581] = 12'b001101110010;
        mem[8582] = 12'b001101110001;
        mem[8583] = 12'b001101110000;
        mem[8584] = 12'b001101110000;
        mem[8585] = 12'b001101101111;
        mem[8586] = 12'b001101101111;
        mem[8587] = 12'b001101101110;
        mem[8588] = 12'b001101101110;
        mem[8589] = 12'b001101101101;
        mem[8590] = 12'b001101101100;
        mem[8591] = 12'b001101101100;
        mem[8592] = 12'b001101101011;
        mem[8593] = 12'b001101101011;
        mem[8594] = 12'b001101101010;
        mem[8595] = 12'b001101101001;
        mem[8596] = 12'b001101101001;
        mem[8597] = 12'b001101101000;
        mem[8598] = 12'b001101101000;
        mem[8599] = 12'b001101100111;
        mem[8600] = 12'b001101100111;
        mem[8601] = 12'b001101100110;
        mem[8602] = 12'b001101100101;
        mem[8603] = 12'b001101100101;
        mem[8604] = 12'b001101100100;
        mem[8605] = 12'b001101100100;
        mem[8606] = 12'b001101100011;
        mem[8607] = 12'b001101100010;
        mem[8608] = 12'b001101100010;
        mem[8609] = 12'b001101100001;
        mem[8610] = 12'b001101100001;
        mem[8611] = 12'b001101100000;
        mem[8612] = 12'b001101100000;
        mem[8613] = 12'b001101011111;
        mem[8614] = 12'b001101011110;
        mem[8615] = 12'b001101011110;
        mem[8616] = 12'b001101011101;
        mem[8617] = 12'b001101011101;
        mem[8618] = 12'b001101011100;
        mem[8619] = 12'b001101011011;
        mem[8620] = 12'b001101011011;
        mem[8621] = 12'b001101011010;
        mem[8622] = 12'b001101011010;
        mem[8623] = 12'b001101011001;
        mem[8624] = 12'b001101011001;
        mem[8625] = 12'b001101011000;
        mem[8626] = 12'b001101010111;
        mem[8627] = 12'b001101010111;
        mem[8628] = 12'b001101010110;
        mem[8629] = 12'b001101010110;
        mem[8630] = 12'b001101010101;
        mem[8631] = 12'b001101010100;
        mem[8632] = 12'b001101010100;
        mem[8633] = 12'b001101010011;
        mem[8634] = 12'b001101010011;
        mem[8635] = 12'b001101010010;
        mem[8636] = 12'b001101010010;
        mem[8637] = 12'b001101010001;
        mem[8638] = 12'b001101010000;
        mem[8639] = 12'b001101010000;
        mem[8640] = 12'b001101001111;
        mem[8641] = 12'b001101001111;
        mem[8642] = 12'b001101001110;
        mem[8643] = 12'b001101001101;
        mem[8644] = 12'b001101001101;
        mem[8645] = 12'b001101001100;
        mem[8646] = 12'b001101001100;
        mem[8647] = 12'b001101001011;
        mem[8648] = 12'b001101001011;
        mem[8649] = 12'b001101001010;
        mem[8650] = 12'b001101001001;
        mem[8651] = 12'b001101001001;
        mem[8652] = 12'b001101001000;
        mem[8653] = 12'b001101001000;
        mem[8654] = 12'b001101000111;
        mem[8655] = 12'b001101000110;
        mem[8656] = 12'b001101000110;
        mem[8657] = 12'b001101000101;
        mem[8658] = 12'b001101000101;
        mem[8659] = 12'b001101000100;
        mem[8660] = 12'b001101000011;
        mem[8661] = 12'b001101000011;
        mem[8662] = 12'b001101000010;
        mem[8663] = 12'b001101000010;
        mem[8664] = 12'b001101000001;
        mem[8665] = 12'b001101000001;
        mem[8666] = 12'b001101000000;
        mem[8667] = 12'b001100111111;
        mem[8668] = 12'b001100111111;
        mem[8669] = 12'b001100111110;
        mem[8670] = 12'b001100111110;
        mem[8671] = 12'b001100111101;
        mem[8672] = 12'b001100111100;
        mem[8673] = 12'b001100111100;
        mem[8674] = 12'b001100111011;
        mem[8675] = 12'b001100111011;
        mem[8676] = 12'b001100111010;
        mem[8677] = 12'b001100111010;
        mem[8678] = 12'b001100111001;
        mem[8679] = 12'b001100111000;
        mem[8680] = 12'b001100111000;
        mem[8681] = 12'b001100110111;
        mem[8682] = 12'b001100110111;
        mem[8683] = 12'b001100110110;
        mem[8684] = 12'b001100110101;
        mem[8685] = 12'b001100110101;
        mem[8686] = 12'b001100110100;
        mem[8687] = 12'b001100110100;
        mem[8688] = 12'b001100110011;
        mem[8689] = 12'b001100110010;
        mem[8690] = 12'b001100110010;
        mem[8691] = 12'b001100110001;
        mem[8692] = 12'b001100110001;
        mem[8693] = 12'b001100110000;
        mem[8694] = 12'b001100101111;
        mem[8695] = 12'b001100101111;
        mem[8696] = 12'b001100101110;
        mem[8697] = 12'b001100101110;
        mem[8698] = 12'b001100101101;
        mem[8699] = 12'b001100101101;
        mem[8700] = 12'b001100101100;
        mem[8701] = 12'b001100101011;
        mem[8702] = 12'b001100101011;
        mem[8703] = 12'b001100101010;
        mem[8704] = 12'b001100101010;
        mem[8705] = 12'b001100101001;
        mem[8706] = 12'b001100101000;
        mem[8707] = 12'b001100101000;
        mem[8708] = 12'b001100100111;
        mem[8709] = 12'b001100100111;
        mem[8710] = 12'b001100100110;
        mem[8711] = 12'b001100100101;
        mem[8712] = 12'b001100100101;
        mem[8713] = 12'b001100100100;
        mem[8714] = 12'b001100100100;
        mem[8715] = 12'b001100100011;
        mem[8716] = 12'b001100100010;
        mem[8717] = 12'b001100100010;
        mem[8718] = 12'b001100100001;
        mem[8719] = 12'b001100100001;
        mem[8720] = 12'b001100100000;
        mem[8721] = 12'b001100100000;
        mem[8722] = 12'b001100011111;
        mem[8723] = 12'b001100011110;
        mem[8724] = 12'b001100011110;
        mem[8725] = 12'b001100011101;
        mem[8726] = 12'b001100011101;
        mem[8727] = 12'b001100011100;
        mem[8728] = 12'b001100011011;
        mem[8729] = 12'b001100011011;
        mem[8730] = 12'b001100011010;
        mem[8731] = 12'b001100011010;
        mem[8732] = 12'b001100011001;
        mem[8733] = 12'b001100011000;
        mem[8734] = 12'b001100011000;
        mem[8735] = 12'b001100010111;
        mem[8736] = 12'b001100010111;
        mem[8737] = 12'b001100010110;
        mem[8738] = 12'b001100010101;
        mem[8739] = 12'b001100010101;
        mem[8740] = 12'b001100010100;
        mem[8741] = 12'b001100010100;
        mem[8742] = 12'b001100010011;
        mem[8743] = 12'b001100010010;
        mem[8744] = 12'b001100010010;
        mem[8745] = 12'b001100010001;
        mem[8746] = 12'b001100010001;
        mem[8747] = 12'b001100010000;
        mem[8748] = 12'b001100010000;
        mem[8749] = 12'b001100001111;
        mem[8750] = 12'b001100001110;
        mem[8751] = 12'b001100001110;
        mem[8752] = 12'b001100001101;
        mem[8753] = 12'b001100001101;
        mem[8754] = 12'b001100001100;
        mem[8755] = 12'b001100001011;
        mem[8756] = 12'b001100001011;
        mem[8757] = 12'b001100001010;
        mem[8758] = 12'b001100001010;
        mem[8759] = 12'b001100001001;
        mem[8760] = 12'b001100001000;
        mem[8761] = 12'b001100001000;
        mem[8762] = 12'b001100000111;
        mem[8763] = 12'b001100000111;
        mem[8764] = 12'b001100000110;
        mem[8765] = 12'b001100000101;
        mem[8766] = 12'b001100000101;
        mem[8767] = 12'b001100000100;
        mem[8768] = 12'b001100000100;
        mem[8769] = 12'b001100000011;
        mem[8770] = 12'b001100000010;
        mem[8771] = 12'b001100000010;
        mem[8772] = 12'b001100000001;
        mem[8773] = 12'b001100000001;
        mem[8774] = 12'b001100000000;
        mem[8775] = 12'b001011111111;
        mem[8776] = 12'b001011111111;
        mem[8777] = 12'b001011111110;
        mem[8778] = 12'b001011111110;
        mem[8779] = 12'b001011111101;
        mem[8780] = 12'b001011111100;
        mem[8781] = 12'b001011111100;
        mem[8782] = 12'b001011111011;
        mem[8783] = 12'b001011111011;
        mem[8784] = 12'b001011111010;
        mem[8785] = 12'b001011111001;
        mem[8786] = 12'b001011111001;
        mem[8787] = 12'b001011111000;
        mem[8788] = 12'b001011111000;
        mem[8789] = 12'b001011110111;
        mem[8790] = 12'b001011110111;
        mem[8791] = 12'b001011110110;
        mem[8792] = 12'b001011110101;
        mem[8793] = 12'b001011110101;
        mem[8794] = 12'b001011110100;
        mem[8795] = 12'b001011110100;
        mem[8796] = 12'b001011110011;
        mem[8797] = 12'b001011110010;
        mem[8798] = 12'b001011110010;
        mem[8799] = 12'b001011110001;
        mem[8800] = 12'b001011110001;
        mem[8801] = 12'b001011110000;
        mem[8802] = 12'b001011101111;
        mem[8803] = 12'b001011101111;
        mem[8804] = 12'b001011101110;
        mem[8805] = 12'b001011101110;
        mem[8806] = 12'b001011101101;
        mem[8807] = 12'b001011101100;
        mem[8808] = 12'b001011101100;
        mem[8809] = 12'b001011101011;
        mem[8810] = 12'b001011101011;
        mem[8811] = 12'b001011101010;
        mem[8812] = 12'b001011101001;
        mem[8813] = 12'b001011101001;
        mem[8814] = 12'b001011101000;
        mem[8815] = 12'b001011101000;
        mem[8816] = 12'b001011100111;
        mem[8817] = 12'b001011100110;
        mem[8818] = 12'b001011100110;
        mem[8819] = 12'b001011100101;
        mem[8820] = 12'b001011100101;
        mem[8821] = 12'b001011100100;
        mem[8822] = 12'b001011100011;
        mem[8823] = 12'b001011100011;
        mem[8824] = 12'b001011100010;
        mem[8825] = 12'b001011100010;
        mem[8826] = 12'b001011100001;
        mem[8827] = 12'b001011100000;
        mem[8828] = 12'b001011100000;
        mem[8829] = 12'b001011011111;
        mem[8830] = 12'b001011011111;
        mem[8831] = 12'b001011011110;
        mem[8832] = 12'b001011011101;
        mem[8833] = 12'b001011011101;
        mem[8834] = 12'b001011011100;
        mem[8835] = 12'b001011011100;
        mem[8836] = 12'b001011011011;
        mem[8837] = 12'b001011011010;
        mem[8838] = 12'b001011011010;
        mem[8839] = 12'b001011011001;
        mem[8840] = 12'b001011011001;
        mem[8841] = 12'b001011011000;
        mem[8842] = 12'b001011010111;
        mem[8843] = 12'b001011010111;
        mem[8844] = 12'b001011010110;
        mem[8845] = 12'b001011010110;
        mem[8846] = 12'b001011010101;
        mem[8847] = 12'b001011010100;
        mem[8848] = 12'b001011010100;
        mem[8849] = 12'b001011010011;
        mem[8850] = 12'b001011010011;
        mem[8851] = 12'b001011010010;
        mem[8852] = 12'b001011010001;
        mem[8853] = 12'b001011010001;
        mem[8854] = 12'b001011010000;
        mem[8855] = 12'b001011010000;
        mem[8856] = 12'b001011001111;
        mem[8857] = 12'b001011001110;
        mem[8858] = 12'b001011001110;
        mem[8859] = 12'b001011001101;
        mem[8860] = 12'b001011001101;
        mem[8861] = 12'b001011001100;
        mem[8862] = 12'b001011001011;
        mem[8863] = 12'b001011001011;
        mem[8864] = 12'b001011001010;
        mem[8865] = 12'b001011001001;
        mem[8866] = 12'b001011001001;
        mem[8867] = 12'b001011001000;
        mem[8868] = 12'b001011001000;
        mem[8869] = 12'b001011000111;
        mem[8870] = 12'b001011000110;
        mem[8871] = 12'b001011000110;
        mem[8872] = 12'b001011000101;
        mem[8873] = 12'b001011000101;
        mem[8874] = 12'b001011000100;
        mem[8875] = 12'b001011000011;
        mem[8876] = 12'b001011000011;
        mem[8877] = 12'b001011000010;
        mem[8878] = 12'b001011000010;
        mem[8879] = 12'b001011000001;
        mem[8880] = 12'b001011000000;
        mem[8881] = 12'b001011000000;
        mem[8882] = 12'b001010111111;
        mem[8883] = 12'b001010111111;
        mem[8884] = 12'b001010111110;
        mem[8885] = 12'b001010111101;
        mem[8886] = 12'b001010111101;
        mem[8887] = 12'b001010111100;
        mem[8888] = 12'b001010111100;
        mem[8889] = 12'b001010111011;
        mem[8890] = 12'b001010111010;
        mem[8891] = 12'b001010111010;
        mem[8892] = 12'b001010111001;
        mem[8893] = 12'b001010111001;
        mem[8894] = 12'b001010111000;
        mem[8895] = 12'b001010110111;
        mem[8896] = 12'b001010110111;
        mem[8897] = 12'b001010110110;
        mem[8898] = 12'b001010110110;
        mem[8899] = 12'b001010110101;
        mem[8900] = 12'b001010110100;
        mem[8901] = 12'b001010110100;
        mem[8902] = 12'b001010110011;
        mem[8903] = 12'b001010110011;
        mem[8904] = 12'b001010110010;
        mem[8905] = 12'b001010110001;
        mem[8906] = 12'b001010110001;
        mem[8907] = 12'b001010110000;
        mem[8908] = 12'b001010110000;
        mem[8909] = 12'b001010101111;
        mem[8910] = 12'b001010101110;
        mem[8911] = 12'b001010101110;
        mem[8912] = 12'b001010101101;
        mem[8913] = 12'b001010101100;
        mem[8914] = 12'b001010101100;
        mem[8915] = 12'b001010101011;
        mem[8916] = 12'b001010101011;
        mem[8917] = 12'b001010101010;
        mem[8918] = 12'b001010101001;
        mem[8919] = 12'b001010101001;
        mem[8920] = 12'b001010101000;
        mem[8921] = 12'b001010101000;
        mem[8922] = 12'b001010100111;
        mem[8923] = 12'b001010100110;
        mem[8924] = 12'b001010100110;
        mem[8925] = 12'b001010100101;
        mem[8926] = 12'b001010100101;
        mem[8927] = 12'b001010100100;
        mem[8928] = 12'b001010100011;
        mem[8929] = 12'b001010100011;
        mem[8930] = 12'b001010100010;
        mem[8931] = 12'b001010100010;
        mem[8932] = 12'b001010100001;
        mem[8933] = 12'b001010100000;
        mem[8934] = 12'b001010100000;
        mem[8935] = 12'b001010011111;
        mem[8936] = 12'b001010011111;
        mem[8937] = 12'b001010011110;
        mem[8938] = 12'b001010011101;
        mem[8939] = 12'b001010011101;
        mem[8940] = 12'b001010011100;
        mem[8941] = 12'b001010011011;
        mem[8942] = 12'b001010011011;
        mem[8943] = 12'b001010011010;
        mem[8944] = 12'b001010011010;
        mem[8945] = 12'b001010011001;
        mem[8946] = 12'b001010011000;
        mem[8947] = 12'b001010011000;
        mem[8948] = 12'b001010010111;
        mem[8949] = 12'b001010010111;
        mem[8950] = 12'b001010010110;
        mem[8951] = 12'b001010010101;
        mem[8952] = 12'b001010010101;
        mem[8953] = 12'b001010010100;
        mem[8954] = 12'b001010010100;
        mem[8955] = 12'b001010010011;
        mem[8956] = 12'b001010010010;
        mem[8957] = 12'b001010010010;
        mem[8958] = 12'b001010010001;
        mem[8959] = 12'b001010010001;
        mem[8960] = 12'b001010010000;
        mem[8961] = 12'b001010001111;
        mem[8962] = 12'b001010001111;
        mem[8963] = 12'b001010001110;
        mem[8964] = 12'b001010001101;
        mem[8965] = 12'b001010001101;
        mem[8966] = 12'b001010001100;
        mem[8967] = 12'b001010001100;
        mem[8968] = 12'b001010001011;
        mem[8969] = 12'b001010001010;
        mem[8970] = 12'b001010001010;
        mem[8971] = 12'b001010001001;
        mem[8972] = 12'b001010001001;
        mem[8973] = 12'b001010001000;
        mem[8974] = 12'b001010000111;
        mem[8975] = 12'b001010000111;
        mem[8976] = 12'b001010000110;
        mem[8977] = 12'b001010000110;
        mem[8978] = 12'b001010000101;
        mem[8979] = 12'b001010000100;
        mem[8980] = 12'b001010000100;
        mem[8981] = 12'b001010000011;
        mem[8982] = 12'b001010000011;
        mem[8983] = 12'b001010000010;
        mem[8984] = 12'b001010000001;
        mem[8985] = 12'b001010000001;
        mem[8986] = 12'b001010000000;
        mem[8987] = 12'b001001111111;
        mem[8988] = 12'b001001111111;
        mem[8989] = 12'b001001111110;
        mem[8990] = 12'b001001111110;
        mem[8991] = 12'b001001111101;
        mem[8992] = 12'b001001111100;
        mem[8993] = 12'b001001111100;
        mem[8994] = 12'b001001111011;
        mem[8995] = 12'b001001111011;
        mem[8996] = 12'b001001111010;
        mem[8997] = 12'b001001111001;
        mem[8998] = 12'b001001111001;
        mem[8999] = 12'b001001111000;
        mem[9000] = 12'b001001111000;
        mem[9001] = 12'b001001110111;
        mem[9002] = 12'b001001110110;
        mem[9003] = 12'b001001110110;
        mem[9004] = 12'b001001110101;
        mem[9005] = 12'b001001110100;
        mem[9006] = 12'b001001110100;
        mem[9007] = 12'b001001110011;
        mem[9008] = 12'b001001110011;
        mem[9009] = 12'b001001110010;
        mem[9010] = 12'b001001110001;
        mem[9011] = 12'b001001110001;
        mem[9012] = 12'b001001110000;
        mem[9013] = 12'b001001110000;
        mem[9014] = 12'b001001101111;
        mem[9015] = 12'b001001101110;
        mem[9016] = 12'b001001101110;
        mem[9017] = 12'b001001101101;
        mem[9018] = 12'b001001101100;
        mem[9019] = 12'b001001101100;
        mem[9020] = 12'b001001101011;
        mem[9021] = 12'b001001101011;
        mem[9022] = 12'b001001101010;
        mem[9023] = 12'b001001101001;
        mem[9024] = 12'b001001101001;
        mem[9025] = 12'b001001101000;
        mem[9026] = 12'b001001101000;
        mem[9027] = 12'b001001100111;
        mem[9028] = 12'b001001100110;
        mem[9029] = 12'b001001100110;
        mem[9030] = 12'b001001100101;
        mem[9031] = 12'b001001100101;
        mem[9032] = 12'b001001100100;
        mem[9033] = 12'b001001100011;
        mem[9034] = 12'b001001100011;
        mem[9035] = 12'b001001100010;
        mem[9036] = 12'b001001100001;
        mem[9037] = 12'b001001100001;
        mem[9038] = 12'b001001100000;
        mem[9039] = 12'b001001100000;
        mem[9040] = 12'b001001011111;
        mem[9041] = 12'b001001011110;
        mem[9042] = 12'b001001011110;
        mem[9043] = 12'b001001011101;
        mem[9044] = 12'b001001011101;
        mem[9045] = 12'b001001011100;
        mem[9046] = 12'b001001011011;
        mem[9047] = 12'b001001011011;
        mem[9048] = 12'b001001011010;
        mem[9049] = 12'b001001011001;
        mem[9050] = 12'b001001011001;
        mem[9051] = 12'b001001011000;
        mem[9052] = 12'b001001011000;
        mem[9053] = 12'b001001010111;
        mem[9054] = 12'b001001010110;
        mem[9055] = 12'b001001010110;
        mem[9056] = 12'b001001010101;
        mem[9057] = 12'b001001010101;
        mem[9058] = 12'b001001010100;
        mem[9059] = 12'b001001010011;
        mem[9060] = 12'b001001010011;
        mem[9061] = 12'b001001010010;
        mem[9062] = 12'b001001010001;
        mem[9063] = 12'b001001010001;
        mem[9064] = 12'b001001010000;
        mem[9065] = 12'b001001010000;
        mem[9066] = 12'b001001001111;
        mem[9067] = 12'b001001001110;
        mem[9068] = 12'b001001001110;
        mem[9069] = 12'b001001001101;
        mem[9070] = 12'b001001001101;
        mem[9071] = 12'b001001001100;
        mem[9072] = 12'b001001001011;
        mem[9073] = 12'b001001001011;
        mem[9074] = 12'b001001001010;
        mem[9075] = 12'b001001001001;
        mem[9076] = 12'b001001001001;
        mem[9077] = 12'b001001001000;
        mem[9078] = 12'b001001001000;
        mem[9079] = 12'b001001000111;
        mem[9080] = 12'b001001000110;
        mem[9081] = 12'b001001000110;
        mem[9082] = 12'b001001000101;
        mem[9083] = 12'b001001000101;
        mem[9084] = 12'b001001000100;
        mem[9085] = 12'b001001000011;
        mem[9086] = 12'b001001000011;
        mem[9087] = 12'b001001000010;
        mem[9088] = 12'b001001000001;
        mem[9089] = 12'b001001000001;
        mem[9090] = 12'b001001000000;
        mem[9091] = 12'b001001000000;
        mem[9092] = 12'b001000111111;
        mem[9093] = 12'b001000111110;
        mem[9094] = 12'b001000111110;
        mem[9095] = 12'b001000111101;
        mem[9096] = 12'b001000111101;
        mem[9097] = 12'b001000111100;
        mem[9098] = 12'b001000111011;
        mem[9099] = 12'b001000111011;
        mem[9100] = 12'b001000111010;
        mem[9101] = 12'b001000111001;
        mem[9102] = 12'b001000111001;
        mem[9103] = 12'b001000111000;
        mem[9104] = 12'b001000111000;
        mem[9105] = 12'b001000110111;
        mem[9106] = 12'b001000110110;
        mem[9107] = 12'b001000110110;
        mem[9108] = 12'b001000110101;
        mem[9109] = 12'b001000110100;
        mem[9110] = 12'b001000110100;
        mem[9111] = 12'b001000110011;
        mem[9112] = 12'b001000110011;
        mem[9113] = 12'b001000110010;
        mem[9114] = 12'b001000110001;
        mem[9115] = 12'b001000110001;
        mem[9116] = 12'b001000110000;
        mem[9117] = 12'b001000110000;
        mem[9118] = 12'b001000101111;
        mem[9119] = 12'b001000101110;
        mem[9120] = 12'b001000101110;
        mem[9121] = 12'b001000101101;
        mem[9122] = 12'b001000101100;
        mem[9123] = 12'b001000101100;
        mem[9124] = 12'b001000101011;
        mem[9125] = 12'b001000101011;
        mem[9126] = 12'b001000101010;
        mem[9127] = 12'b001000101001;
        mem[9128] = 12'b001000101001;
        mem[9129] = 12'b001000101000;
        mem[9130] = 12'b001000100111;
        mem[9131] = 12'b001000100111;
        mem[9132] = 12'b001000100110;
        mem[9133] = 12'b001000100110;
        mem[9134] = 12'b001000100101;
        mem[9135] = 12'b001000100100;
        mem[9136] = 12'b001000100100;
        mem[9137] = 12'b001000100011;
        mem[9138] = 12'b001000100011;
        mem[9139] = 12'b001000100010;
        mem[9140] = 12'b001000100001;
        mem[9141] = 12'b001000100001;
        mem[9142] = 12'b001000100000;
        mem[9143] = 12'b001000011111;
        mem[9144] = 12'b001000011111;
        mem[9145] = 12'b001000011110;
        mem[9146] = 12'b001000011110;
        mem[9147] = 12'b001000011101;
        mem[9148] = 12'b001000011100;
        mem[9149] = 12'b001000011100;
        mem[9150] = 12'b001000011011;
        mem[9151] = 12'b001000011010;
        mem[9152] = 12'b001000011010;
        mem[9153] = 12'b001000011001;
        mem[9154] = 12'b001000011001;
        mem[9155] = 12'b001000011000;
        mem[9156] = 12'b001000010111;
        mem[9157] = 12'b001000010111;
        mem[9158] = 12'b001000010110;
        mem[9159] = 12'b001000010101;
        mem[9160] = 12'b001000010101;
        mem[9161] = 12'b001000010100;
        mem[9162] = 12'b001000010100;
        mem[9163] = 12'b001000010011;
        mem[9164] = 12'b001000010010;
        mem[9165] = 12'b001000010010;
        mem[9166] = 12'b001000010001;
        mem[9167] = 12'b001000010001;
        mem[9168] = 12'b001000010000;
        mem[9169] = 12'b001000001111;
        mem[9170] = 12'b001000001111;
        mem[9171] = 12'b001000001110;
        mem[9172] = 12'b001000001101;
        mem[9173] = 12'b001000001101;
        mem[9174] = 12'b001000001100;
        mem[9175] = 12'b001000001100;
        mem[9176] = 12'b001000001011;
        mem[9177] = 12'b001000001010;
        mem[9178] = 12'b001000001010;
        mem[9179] = 12'b001000001001;
        mem[9180] = 12'b001000001000;
        mem[9181] = 12'b001000001000;
        mem[9182] = 12'b001000000111;
        mem[9183] = 12'b001000000111;
        mem[9184] = 12'b001000000110;
        mem[9185] = 12'b001000000101;
        mem[9186] = 12'b001000000101;
        mem[9187] = 12'b001000000100;
        mem[9188] = 12'b001000000011;
        mem[9189] = 12'b001000000011;
        mem[9190] = 12'b001000000010;
        mem[9191] = 12'b001000000010;
        mem[9192] = 12'b001000000001;
        mem[9193] = 12'b001000000000;
        mem[9194] = 12'b001000000000;
        mem[9195] = 12'b000111111111;
        mem[9196] = 12'b000111111110;
        mem[9197] = 12'b000111111110;
        mem[9198] = 12'b000111111101;
        mem[9199] = 12'b000111111101;
        mem[9200] = 12'b000111111100;
        mem[9201] = 12'b000111111011;
        mem[9202] = 12'b000111111011;
        mem[9203] = 12'b000111111010;
        mem[9204] = 12'b000111111010;
        mem[9205] = 12'b000111111001;
        mem[9206] = 12'b000111111000;
        mem[9207] = 12'b000111111000;
        mem[9208] = 12'b000111110111;
        mem[9209] = 12'b000111110110;
        mem[9210] = 12'b000111110110;
        mem[9211] = 12'b000111110101;
        mem[9212] = 12'b000111110101;
        mem[9213] = 12'b000111110100;
        mem[9214] = 12'b000111110011;
        mem[9215] = 12'b000111110011;
        mem[9216] = 12'b000111110010;
        mem[9217] = 12'b000111110001;
        mem[9218] = 12'b000111110001;
        mem[9219] = 12'b000111110000;
        mem[9220] = 12'b000111110000;
        mem[9221] = 12'b000111101111;
        mem[9222] = 12'b000111101110;
        mem[9223] = 12'b000111101110;
        mem[9224] = 12'b000111101101;
        mem[9225] = 12'b000111101100;
        mem[9226] = 12'b000111101100;
        mem[9227] = 12'b000111101011;
        mem[9228] = 12'b000111101011;
        mem[9229] = 12'b000111101010;
        mem[9230] = 12'b000111101001;
        mem[9231] = 12'b000111101001;
        mem[9232] = 12'b000111101000;
        mem[9233] = 12'b000111100111;
        mem[9234] = 12'b000111100111;
        mem[9235] = 12'b000111100110;
        mem[9236] = 12'b000111100110;
        mem[9237] = 12'b000111100101;
        mem[9238] = 12'b000111100100;
        mem[9239] = 12'b000111100100;
        mem[9240] = 12'b000111100011;
        mem[9241] = 12'b000111100010;
        mem[9242] = 12'b000111100010;
        mem[9243] = 12'b000111100001;
        mem[9244] = 12'b000111100001;
        mem[9245] = 12'b000111100000;
        mem[9246] = 12'b000111011111;
        mem[9247] = 12'b000111011111;
        mem[9248] = 12'b000111011110;
        mem[9249] = 12'b000111011101;
        mem[9250] = 12'b000111011101;
        mem[9251] = 12'b000111011100;
        mem[9252] = 12'b000111011100;
        mem[9253] = 12'b000111011011;
        mem[9254] = 12'b000111011010;
        mem[9255] = 12'b000111011010;
        mem[9256] = 12'b000111011001;
        mem[9257] = 12'b000111011000;
        mem[9258] = 12'b000111011000;
        mem[9259] = 12'b000111010111;
        mem[9260] = 12'b000111010111;
        mem[9261] = 12'b000111010110;
        mem[9262] = 12'b000111010101;
        mem[9263] = 12'b000111010101;
        mem[9264] = 12'b000111010100;
        mem[9265] = 12'b000111010011;
        mem[9266] = 12'b000111010011;
        mem[9267] = 12'b000111010010;
        mem[9268] = 12'b000111010010;
        mem[9269] = 12'b000111010001;
        mem[9270] = 12'b000111010000;
        mem[9271] = 12'b000111010000;
        mem[9272] = 12'b000111001111;
        mem[9273] = 12'b000111001110;
        mem[9274] = 12'b000111001110;
        mem[9275] = 12'b000111001101;
        mem[9276] = 12'b000111001101;
        mem[9277] = 12'b000111001100;
        mem[9278] = 12'b000111001011;
        mem[9279] = 12'b000111001011;
        mem[9280] = 12'b000111001010;
        mem[9281] = 12'b000111001001;
        mem[9282] = 12'b000111001001;
        mem[9283] = 12'b000111001000;
        mem[9284] = 12'b000111000111;
        mem[9285] = 12'b000111000111;
        mem[9286] = 12'b000111000110;
        mem[9287] = 12'b000111000110;
        mem[9288] = 12'b000111000101;
        mem[9289] = 12'b000111000100;
        mem[9290] = 12'b000111000100;
        mem[9291] = 12'b000111000011;
        mem[9292] = 12'b000111000010;
        mem[9293] = 12'b000111000010;
        mem[9294] = 12'b000111000001;
        mem[9295] = 12'b000111000001;
        mem[9296] = 12'b000111000000;
        mem[9297] = 12'b000110111111;
        mem[9298] = 12'b000110111111;
        mem[9299] = 12'b000110111110;
        mem[9300] = 12'b000110111101;
        mem[9301] = 12'b000110111101;
        mem[9302] = 12'b000110111100;
        mem[9303] = 12'b000110111100;
        mem[9304] = 12'b000110111011;
        mem[9305] = 12'b000110111010;
        mem[9306] = 12'b000110111010;
        mem[9307] = 12'b000110111001;
        mem[9308] = 12'b000110111000;
        mem[9309] = 12'b000110111000;
        mem[9310] = 12'b000110110111;
        mem[9311] = 12'b000110110111;
        mem[9312] = 12'b000110110110;
        mem[9313] = 12'b000110110101;
        mem[9314] = 12'b000110110101;
        mem[9315] = 12'b000110110100;
        mem[9316] = 12'b000110110011;
        mem[9317] = 12'b000110110011;
        mem[9318] = 12'b000110110010;
        mem[9319] = 12'b000110110010;
        mem[9320] = 12'b000110110001;
        mem[9321] = 12'b000110110000;
        mem[9322] = 12'b000110110000;
        mem[9323] = 12'b000110101111;
        mem[9324] = 12'b000110101110;
        mem[9325] = 12'b000110101110;
        mem[9326] = 12'b000110101101;
        mem[9327] = 12'b000110101100;
        mem[9328] = 12'b000110101100;
        mem[9329] = 12'b000110101011;
        mem[9330] = 12'b000110101011;
        mem[9331] = 12'b000110101010;
        mem[9332] = 12'b000110101001;
        mem[9333] = 12'b000110101001;
        mem[9334] = 12'b000110101000;
        mem[9335] = 12'b000110100111;
        mem[9336] = 12'b000110100111;
        mem[9337] = 12'b000110100110;
        mem[9338] = 12'b000110100110;
        mem[9339] = 12'b000110100101;
        mem[9340] = 12'b000110100100;
        mem[9341] = 12'b000110100100;
        mem[9342] = 12'b000110100011;
        mem[9343] = 12'b000110100010;
        mem[9344] = 12'b000110100010;
        mem[9345] = 12'b000110100001;
        mem[9346] = 12'b000110100001;
        mem[9347] = 12'b000110100000;
        mem[9348] = 12'b000110011111;
        mem[9349] = 12'b000110011111;
        mem[9350] = 12'b000110011110;
        mem[9351] = 12'b000110011101;
        mem[9352] = 12'b000110011101;
        mem[9353] = 12'b000110011100;
        mem[9354] = 12'b000110011011;
        mem[9355] = 12'b000110011011;
        mem[9356] = 12'b000110011010;
        mem[9357] = 12'b000110011010;
        mem[9358] = 12'b000110011001;
        mem[9359] = 12'b000110011000;
        mem[9360] = 12'b000110011000;
        mem[9361] = 12'b000110010111;
        mem[9362] = 12'b000110010110;
        mem[9363] = 12'b000110010110;
        mem[9364] = 12'b000110010101;
        mem[9365] = 12'b000110010101;
        mem[9366] = 12'b000110010100;
        mem[9367] = 12'b000110010011;
        mem[9368] = 12'b000110010011;
        mem[9369] = 12'b000110010010;
        mem[9370] = 12'b000110010001;
        mem[9371] = 12'b000110010001;
        mem[9372] = 12'b000110010000;
        mem[9373] = 12'b000110010000;
        mem[9374] = 12'b000110001111;
        mem[9375] = 12'b000110001110;
        mem[9376] = 12'b000110001110;
        mem[9377] = 12'b000110001101;
        mem[9378] = 12'b000110001100;
        mem[9379] = 12'b000110001100;
        mem[9380] = 12'b000110001011;
        mem[9381] = 12'b000110001010;
        mem[9382] = 12'b000110001010;
        mem[9383] = 12'b000110001001;
        mem[9384] = 12'b000110001001;
        mem[9385] = 12'b000110001000;
        mem[9386] = 12'b000110000111;
        mem[9387] = 12'b000110000111;
        mem[9388] = 12'b000110000110;
        mem[9389] = 12'b000110000101;
        mem[9390] = 12'b000110000101;
        mem[9391] = 12'b000110000100;
        mem[9392] = 12'b000110000100;
        mem[9393] = 12'b000110000011;
        mem[9394] = 12'b000110000010;
        mem[9395] = 12'b000110000010;
        mem[9396] = 12'b000110000001;
        mem[9397] = 12'b000110000000;
        mem[9398] = 12'b000110000000;
        mem[9399] = 12'b000101111111;
        mem[9400] = 12'b000101111110;
        mem[9401] = 12'b000101111110;
        mem[9402] = 12'b000101111101;
        mem[9403] = 12'b000101111101;
        mem[9404] = 12'b000101111100;
        mem[9405] = 12'b000101111011;
        mem[9406] = 12'b000101111011;
        mem[9407] = 12'b000101111010;
        mem[9408] = 12'b000101111001;
        mem[9409] = 12'b000101111001;
        mem[9410] = 12'b000101111000;
        mem[9411] = 12'b000101111000;
        mem[9412] = 12'b000101110111;
        mem[9413] = 12'b000101110110;
        mem[9414] = 12'b000101110110;
        mem[9415] = 12'b000101110101;
        mem[9416] = 12'b000101110100;
        mem[9417] = 12'b000101110100;
        mem[9418] = 12'b000101110011;
        mem[9419] = 12'b000101110010;
        mem[9420] = 12'b000101110010;
        mem[9421] = 12'b000101110001;
        mem[9422] = 12'b000101110001;
        mem[9423] = 12'b000101110000;
        mem[9424] = 12'b000101101111;
        mem[9425] = 12'b000101101111;
        mem[9426] = 12'b000101101110;
        mem[9427] = 12'b000101101101;
        mem[9428] = 12'b000101101101;
        mem[9429] = 12'b000101101100;
        mem[9430] = 12'b000101101100;
        mem[9431] = 12'b000101101011;
        mem[9432] = 12'b000101101010;
        mem[9433] = 12'b000101101010;
        mem[9434] = 12'b000101101001;
        mem[9435] = 12'b000101101000;
        mem[9436] = 12'b000101101000;
        mem[9437] = 12'b000101100111;
        mem[9438] = 12'b000101100110;
        mem[9439] = 12'b000101100110;
        mem[9440] = 12'b000101100101;
        mem[9441] = 12'b000101100101;
        mem[9442] = 12'b000101100100;
        mem[9443] = 12'b000101100011;
        mem[9444] = 12'b000101100011;
        mem[9445] = 12'b000101100010;
        mem[9446] = 12'b000101100001;
        mem[9447] = 12'b000101100001;
        mem[9448] = 12'b000101100000;
        mem[9449] = 12'b000101011111;
        mem[9450] = 12'b000101011111;
        mem[9451] = 12'b000101011110;
        mem[9452] = 12'b000101011110;
        mem[9453] = 12'b000101011101;
        mem[9454] = 12'b000101011100;
        mem[9455] = 12'b000101011100;
        mem[9456] = 12'b000101011011;
        mem[9457] = 12'b000101011010;
        mem[9458] = 12'b000101011010;
        mem[9459] = 12'b000101011001;
        mem[9460] = 12'b000101011001;
        mem[9461] = 12'b000101011000;
        mem[9462] = 12'b000101010111;
        mem[9463] = 12'b000101010111;
        mem[9464] = 12'b000101010110;
        mem[9465] = 12'b000101010101;
        mem[9466] = 12'b000101010101;
        mem[9467] = 12'b000101010100;
        mem[9468] = 12'b000101010011;
        mem[9469] = 12'b000101010011;
        mem[9470] = 12'b000101010010;
        mem[9471] = 12'b000101010010;
        mem[9472] = 12'b000101010001;
        mem[9473] = 12'b000101010000;
        mem[9474] = 12'b000101010000;
        mem[9475] = 12'b000101001111;
        mem[9476] = 12'b000101001110;
        mem[9477] = 12'b000101001110;
        mem[9478] = 12'b000101001101;
        mem[9479] = 12'b000101001100;
        mem[9480] = 12'b000101001100;
        mem[9481] = 12'b000101001011;
        mem[9482] = 12'b000101001011;
        mem[9483] = 12'b000101001010;
        mem[9484] = 12'b000101001001;
        mem[9485] = 12'b000101001001;
        mem[9486] = 12'b000101001000;
        mem[9487] = 12'b000101000111;
        mem[9488] = 12'b000101000111;
        mem[9489] = 12'b000101000110;
        mem[9490] = 12'b000101000101;
        mem[9491] = 12'b000101000101;
        mem[9492] = 12'b000101000100;
        mem[9493] = 12'b000101000100;
        mem[9494] = 12'b000101000011;
        mem[9495] = 12'b000101000010;
        mem[9496] = 12'b000101000010;
        mem[9497] = 12'b000101000001;
        mem[9498] = 12'b000101000000;
        mem[9499] = 12'b000101000000;
        mem[9500] = 12'b000100111111;
        mem[9501] = 12'b000100111110;
        mem[9502] = 12'b000100111110;
        mem[9503] = 12'b000100111101;
        mem[9504] = 12'b000100111101;
        mem[9505] = 12'b000100111100;
        mem[9506] = 12'b000100111011;
        mem[9507] = 12'b000100111011;
        mem[9508] = 12'b000100111010;
        mem[9509] = 12'b000100111001;
        mem[9510] = 12'b000100111001;
        mem[9511] = 12'b000100111000;
        mem[9512] = 12'b000100110111;
        mem[9513] = 12'b000100110111;
        mem[9514] = 12'b000100110110;
        mem[9515] = 12'b000100110110;
        mem[9516] = 12'b000100110101;
        mem[9517] = 12'b000100110100;
        mem[9518] = 12'b000100110100;
        mem[9519] = 12'b000100110011;
        mem[9520] = 12'b000100110010;
        mem[9521] = 12'b000100110010;
        mem[9522] = 12'b000100110001;
        mem[9523] = 12'b000100110000;
        mem[9524] = 12'b000100110000;
        mem[9525] = 12'b000100101111;
        mem[9526] = 12'b000100101111;
        mem[9527] = 12'b000100101110;
        mem[9528] = 12'b000100101101;
        mem[9529] = 12'b000100101101;
        mem[9530] = 12'b000100101100;
        mem[9531] = 12'b000100101011;
        mem[9532] = 12'b000100101011;
        mem[9533] = 12'b000100101010;
        mem[9534] = 12'b000100101010;
        mem[9535] = 12'b000100101001;
        mem[9536] = 12'b000100101000;
        mem[9537] = 12'b000100101000;
        mem[9538] = 12'b000100100111;
        mem[9539] = 12'b000100100110;
        mem[9540] = 12'b000100100110;
        mem[9541] = 12'b000100100101;
        mem[9542] = 12'b000100100100;
        mem[9543] = 12'b000100100100;
        mem[9544] = 12'b000100100011;
        mem[9545] = 12'b000100100011;
        mem[9546] = 12'b000100100010;
        mem[9547] = 12'b000100100001;
        mem[9548] = 12'b000100100001;
        mem[9549] = 12'b000100100000;
        mem[9550] = 12'b000100011111;
        mem[9551] = 12'b000100011111;
        mem[9552] = 12'b000100011110;
        mem[9553] = 12'b000100011101;
        mem[9554] = 12'b000100011101;
        mem[9555] = 12'b000100011100;
        mem[9556] = 12'b000100011011;
        mem[9557] = 12'b000100011011;
        mem[9558] = 12'b000100011010;
        mem[9559] = 12'b000100011010;
        mem[9560] = 12'b000100011001;
        mem[9561] = 12'b000100011000;
        mem[9562] = 12'b000100011000;
        mem[9563] = 12'b000100010111;
        mem[9564] = 12'b000100010110;
        mem[9565] = 12'b000100010110;
        mem[9566] = 12'b000100010101;
        mem[9567] = 12'b000100010100;
        mem[9568] = 12'b000100010100;
        mem[9569] = 12'b000100010011;
        mem[9570] = 12'b000100010011;
        mem[9571] = 12'b000100010010;
        mem[9572] = 12'b000100010001;
        mem[9573] = 12'b000100010001;
        mem[9574] = 12'b000100010000;
        mem[9575] = 12'b000100001111;
        mem[9576] = 12'b000100001111;
        mem[9577] = 12'b000100001110;
        mem[9578] = 12'b000100001101;
        mem[9579] = 12'b000100001101;
        mem[9580] = 12'b000100001100;
        mem[9581] = 12'b000100001100;
        mem[9582] = 12'b000100001011;
        mem[9583] = 12'b000100001010;
        mem[9584] = 12'b000100001010;
        mem[9585] = 12'b000100001001;
        mem[9586] = 12'b000100001000;
        mem[9587] = 12'b000100001000;
        mem[9588] = 12'b000100000111;
        mem[9589] = 12'b000100000110;
        mem[9590] = 12'b000100000110;
        mem[9591] = 12'b000100000101;
        mem[9592] = 12'b000100000101;
        mem[9593] = 12'b000100000100;
        mem[9594] = 12'b000100000011;
        mem[9595] = 12'b000100000011;
        mem[9596] = 12'b000100000010;
        mem[9597] = 12'b000100000001;
        mem[9598] = 12'b000100000001;
        mem[9599] = 12'b000100000000;
        mem[9600] = 12'b000011111111;
        mem[9601] = 12'b000011111111;
        mem[9602] = 12'b000011111110;
        mem[9603] = 12'b000011111110;
        mem[9604] = 12'b000011111101;
        mem[9605] = 12'b000011111100;
        mem[9606] = 12'b000011111100;
        mem[9607] = 12'b000011111011;
        mem[9608] = 12'b000011111010;
        mem[9609] = 12'b000011111010;
        mem[9610] = 12'b000011111001;
        mem[9611] = 12'b000011111000;
        mem[9612] = 12'b000011111000;
        mem[9613] = 12'b000011110111;
        mem[9614] = 12'b000011110111;
        mem[9615] = 12'b000011110110;
        mem[9616] = 12'b000011110101;
        mem[9617] = 12'b000011110101;
        mem[9618] = 12'b000011110100;
        mem[9619] = 12'b000011110011;
        mem[9620] = 12'b000011110011;
        mem[9621] = 12'b000011110010;
        mem[9622] = 12'b000011110001;
        mem[9623] = 12'b000011110001;
        mem[9624] = 12'b000011110000;
        mem[9625] = 12'b000011101111;
        mem[9626] = 12'b000011101111;
        mem[9627] = 12'b000011101110;
        mem[9628] = 12'b000011101110;
        mem[9629] = 12'b000011101101;
        mem[9630] = 12'b000011101100;
        mem[9631] = 12'b000011101100;
        mem[9632] = 12'b000011101011;
        mem[9633] = 12'b000011101010;
        mem[9634] = 12'b000011101010;
        mem[9635] = 12'b000011101001;
        mem[9636] = 12'b000011101000;
        mem[9637] = 12'b000011101000;
        mem[9638] = 12'b000011100111;
        mem[9639] = 12'b000011100111;
        mem[9640] = 12'b000011100110;
        mem[9641] = 12'b000011100101;
        mem[9642] = 12'b000011100101;
        mem[9643] = 12'b000011100100;
        mem[9644] = 12'b000011100011;
        mem[9645] = 12'b000011100011;
        mem[9646] = 12'b000011100010;
        mem[9647] = 12'b000011100001;
        mem[9648] = 12'b000011100001;
        mem[9649] = 12'b000011100000;
        mem[9650] = 12'b000011100000;
        mem[9651] = 12'b000011011111;
        mem[9652] = 12'b000011011110;
        mem[9653] = 12'b000011011110;
        mem[9654] = 12'b000011011101;
        mem[9655] = 12'b000011011100;
        mem[9656] = 12'b000011011100;
        mem[9657] = 12'b000011011011;
        mem[9658] = 12'b000011011010;
        mem[9659] = 12'b000011011010;
        mem[9660] = 12'b000011011001;
        mem[9661] = 12'b000011011000;
        mem[9662] = 12'b000011011000;
        mem[9663] = 12'b000011010111;
        mem[9664] = 12'b000011010111;
        mem[9665] = 12'b000011010110;
        mem[9666] = 12'b000011010101;
        mem[9667] = 12'b000011010101;
        mem[9668] = 12'b000011010100;
        mem[9669] = 12'b000011010011;
        mem[9670] = 12'b000011010011;
        mem[9671] = 12'b000011010010;
        mem[9672] = 12'b000011010001;
        mem[9673] = 12'b000011010001;
        mem[9674] = 12'b000011010000;
        mem[9675] = 12'b000011010000;
        mem[9676] = 12'b000011001111;
        mem[9677] = 12'b000011001110;
        mem[9678] = 12'b000011001110;
        mem[9679] = 12'b000011001101;
        mem[9680] = 12'b000011001100;
        mem[9681] = 12'b000011001100;
        mem[9682] = 12'b000011001011;
        mem[9683] = 12'b000011001010;
        mem[9684] = 12'b000011001010;
        mem[9685] = 12'b000011001001;
        mem[9686] = 12'b000011001000;
        mem[9687] = 12'b000011001000;
        mem[9688] = 12'b000011000111;
        mem[9689] = 12'b000011000111;
        mem[9690] = 12'b000011000110;
        mem[9691] = 12'b000011000101;
        mem[9692] = 12'b000011000101;
        mem[9693] = 12'b000011000100;
        mem[9694] = 12'b000011000011;
        mem[9695] = 12'b000011000011;
        mem[9696] = 12'b000011000010;
        mem[9697] = 12'b000011000001;
        mem[9698] = 12'b000011000001;
        mem[9699] = 12'b000011000000;
        mem[9700] = 12'b000011000000;
        mem[9701] = 12'b000010111111;
        mem[9702] = 12'b000010111110;
        mem[9703] = 12'b000010111110;
        mem[9704] = 12'b000010111101;
        mem[9705] = 12'b000010111100;
        mem[9706] = 12'b000010111100;
        mem[9707] = 12'b000010111011;
        mem[9708] = 12'b000010111010;
        mem[9709] = 12'b000010111010;
        mem[9710] = 12'b000010111001;
        mem[9711] = 12'b000010111000;
        mem[9712] = 12'b000010111000;
        mem[9713] = 12'b000010110111;
        mem[9714] = 12'b000010110111;
        mem[9715] = 12'b000010110110;
        mem[9716] = 12'b000010110101;
        mem[9717] = 12'b000010110101;
        mem[9718] = 12'b000010110100;
        mem[9719] = 12'b000010110011;
        mem[9720] = 12'b000010110011;
        mem[9721] = 12'b000010110010;
        mem[9722] = 12'b000010110001;
        mem[9723] = 12'b000010110001;
        mem[9724] = 12'b000010110000;
        mem[9725] = 12'b000010110000;
        mem[9726] = 12'b000010101111;
        mem[9727] = 12'b000010101110;
        mem[9728] = 12'b000010101110;
        mem[9729] = 12'b000010101101;
        mem[9730] = 12'b000010101100;
        mem[9731] = 12'b000010101100;
        mem[9732] = 12'b000010101011;
        mem[9733] = 12'b000010101010;
        mem[9734] = 12'b000010101010;
        mem[9735] = 12'b000010101001;
        mem[9736] = 12'b000010101000;
        mem[9737] = 12'b000010101000;
        mem[9738] = 12'b000010100111;
        mem[9739] = 12'b000010100111;
        mem[9740] = 12'b000010100110;
        mem[9741] = 12'b000010100101;
        mem[9742] = 12'b000010100101;
        mem[9743] = 12'b000010100100;
        mem[9744] = 12'b000010100011;
        mem[9745] = 12'b000010100011;
        mem[9746] = 12'b000010100010;
        mem[9747] = 12'b000010100001;
        mem[9748] = 12'b000010100001;
        mem[9749] = 12'b000010100000;
        mem[9750] = 12'b000010011111;
        mem[9751] = 12'b000010011111;
        mem[9752] = 12'b000010011110;
        mem[9753] = 12'b000010011110;
        mem[9754] = 12'b000010011101;
        mem[9755] = 12'b000010011100;
        mem[9756] = 12'b000010011100;
        mem[9757] = 12'b000010011011;
        mem[9758] = 12'b000010011010;
        mem[9759] = 12'b000010011010;
        mem[9760] = 12'b000010011001;
        mem[9761] = 12'b000010011000;
        mem[9762] = 12'b000010011000;
        mem[9763] = 12'b000010010111;
        mem[9764] = 12'b000010010111;
        mem[9765] = 12'b000010010110;
        mem[9766] = 12'b000010010101;
        mem[9767] = 12'b000010010101;
        mem[9768] = 12'b000010010100;
        mem[9769] = 12'b000010010011;
        mem[9770] = 12'b000010010011;
        mem[9771] = 12'b000010010010;
        mem[9772] = 12'b000010010001;
        mem[9773] = 12'b000010010001;
        mem[9774] = 12'b000010010000;
        mem[9775] = 12'b000010001111;
        mem[9776] = 12'b000010001111;
        mem[9777] = 12'b000010001110;
        mem[9778] = 12'b000010001110;
        mem[9779] = 12'b000010001101;
        mem[9780] = 12'b000010001100;
        mem[9781] = 12'b000010001100;
        mem[9782] = 12'b000010001011;
        mem[9783] = 12'b000010001010;
        mem[9784] = 12'b000010001010;
        mem[9785] = 12'b000010001001;
        mem[9786] = 12'b000010001000;
        mem[9787] = 12'b000010001000;
        mem[9788] = 12'b000010000111;
        mem[9789] = 12'b000010000110;
        mem[9790] = 12'b000010000110;
        mem[9791] = 12'b000010000101;
        mem[9792] = 12'b000010000101;
        mem[9793] = 12'b000010000100;
        mem[9794] = 12'b000010000011;
        mem[9795] = 12'b000010000011;
        mem[9796] = 12'b000010000010;
        mem[9797] = 12'b000010000001;
        mem[9798] = 12'b000010000001;
        mem[9799] = 12'b000010000000;
        mem[9800] = 12'b000001111111;
        mem[9801] = 12'b000001111111;
        mem[9802] = 12'b000001111110;
        mem[9803] = 12'b000001111101;
        mem[9804] = 12'b000001111101;
        mem[9805] = 12'b000001111100;
        mem[9806] = 12'b000001111100;
        mem[9807] = 12'b000001111011;
        mem[9808] = 12'b000001111010;
        mem[9809] = 12'b000001111010;
        mem[9810] = 12'b000001111001;
        mem[9811] = 12'b000001111000;
        mem[9812] = 12'b000001111000;
        mem[9813] = 12'b000001110111;
        mem[9814] = 12'b000001110110;
        mem[9815] = 12'b000001110110;
        mem[9816] = 12'b000001110101;
        mem[9817] = 12'b000001110100;
        mem[9818] = 12'b000001110100;
        mem[9819] = 12'b000001110011;
        mem[9820] = 12'b000001110011;
        mem[9821] = 12'b000001110010;
        mem[9822] = 12'b000001110001;
        mem[9823] = 12'b000001110001;
        mem[9824] = 12'b000001110000;
        mem[9825] = 12'b000001101111;
        mem[9826] = 12'b000001101111;
        mem[9827] = 12'b000001101110;
        mem[9828] = 12'b000001101101;
        mem[9829] = 12'b000001101101;
        mem[9830] = 12'b000001101100;
        mem[9831] = 12'b000001101011;
        mem[9832] = 12'b000001101011;
        mem[9833] = 12'b000001101010;
        mem[9834] = 12'b000001101010;
        mem[9835] = 12'b000001101001;
        mem[9836] = 12'b000001101000;
        mem[9837] = 12'b000001101000;
        mem[9838] = 12'b000001100111;
        mem[9839] = 12'b000001100110;
        mem[9840] = 12'b000001100110;
        mem[9841] = 12'b000001100101;
        mem[9842] = 12'b000001100100;
        mem[9843] = 12'b000001100100;
        mem[9844] = 12'b000001100011;
        mem[9845] = 12'b000001100011;
        mem[9846] = 12'b000001100010;
        mem[9847] = 12'b000001100001;
        mem[9848] = 12'b000001100001;
        mem[9849] = 12'b000001100000;
        mem[9850] = 12'b000001011111;
        mem[9851] = 12'b000001011111;
        mem[9852] = 12'b000001011110;
        mem[9853] = 12'b000001011101;
        mem[9854] = 12'b000001011101;
        mem[9855] = 12'b000001011100;
        mem[9856] = 12'b000001011011;
        mem[9857] = 12'b000001011011;
        mem[9858] = 12'b000001011010;
        mem[9859] = 12'b000001011010;
        mem[9860] = 12'b000001011001;
        mem[9861] = 12'b000001011000;
        mem[9862] = 12'b000001011000;
        mem[9863] = 12'b000001010111;
        mem[9864] = 12'b000001010110;
        mem[9865] = 12'b000001010110;
        mem[9866] = 12'b000001010101;
        mem[9867] = 12'b000001010100;
        mem[9868] = 12'b000001010100;
        mem[9869] = 12'b000001010011;
        mem[9870] = 12'b000001010010;
        mem[9871] = 12'b000001010010;
        mem[9872] = 12'b000001010001;
        mem[9873] = 12'b000001010001;
        mem[9874] = 12'b000001010000;
        mem[9875] = 12'b000001001111;
        mem[9876] = 12'b000001001111;
        mem[9877] = 12'b000001001110;
        mem[9878] = 12'b000001001101;
        mem[9879] = 12'b000001001101;
        mem[9880] = 12'b000001001100;
        mem[9881] = 12'b000001001011;
        mem[9882] = 12'b000001001011;
        mem[9883] = 12'b000001001010;
        mem[9884] = 12'b000001001001;
        mem[9885] = 12'b000001001001;
        mem[9886] = 12'b000001001000;
        mem[9887] = 12'b000001001000;
        mem[9888] = 12'b000001000111;
        mem[9889] = 12'b000001000110;
        mem[9890] = 12'b000001000110;
        mem[9891] = 12'b000001000101;
        mem[9892] = 12'b000001000100;
        mem[9893] = 12'b000001000100;
        mem[9894] = 12'b000001000011;
        mem[9895] = 12'b000001000010;
        mem[9896] = 12'b000001000010;
        mem[9897] = 12'b000001000001;
        mem[9898] = 12'b000001000000;
        mem[9899] = 12'b000001000000;
        mem[9900] = 12'b000000111111;
        mem[9901] = 12'b000000111111;
        mem[9902] = 12'b000000111110;
        mem[9903] = 12'b000000111101;
        mem[9904] = 12'b000000111101;
        mem[9905] = 12'b000000111100;
        mem[9906] = 12'b000000111011;
        mem[9907] = 12'b000000111011;
        mem[9908] = 12'b000000111010;
        mem[9909] = 12'b000000111001;
        mem[9910] = 12'b000000111001;
        mem[9911] = 12'b000000111000;
        mem[9912] = 12'b000000110111;
        mem[9913] = 12'b000000110111;
        mem[9914] = 12'b000000110110;
        mem[9915] = 12'b000000110110;
        mem[9916] = 12'b000000110101;
        mem[9917] = 12'b000000110100;
        mem[9918] = 12'b000000110100;
        mem[9919] = 12'b000000110011;
        mem[9920] = 12'b000000110010;
        mem[9921] = 12'b000000110010;
        mem[9922] = 12'b000000110001;
        mem[9923] = 12'b000000110000;
        mem[9924] = 12'b000000110000;
        mem[9925] = 12'b000000101111;
        mem[9926] = 12'b000000101110;
        mem[9927] = 12'b000000101110;
        mem[9928] = 12'b000000101101;
        mem[9929] = 12'b000000101101;
        mem[9930] = 12'b000000101100;
        mem[9931] = 12'b000000101011;
        mem[9932] = 12'b000000101011;
        mem[9933] = 12'b000000101010;
        mem[9934] = 12'b000000101001;
        mem[9935] = 12'b000000101001;
        mem[9936] = 12'b000000101000;
        mem[9937] = 12'b000000100111;
        mem[9938] = 12'b000000100111;
        mem[9939] = 12'b000000100110;
        mem[9940] = 12'b000000100101;
        mem[9941] = 12'b000000100101;
        mem[9942] = 12'b000000100100;
        mem[9943] = 12'b000000100100;
        mem[9944] = 12'b000000100011;
        mem[9945] = 12'b000000100010;
        mem[9946] = 12'b000000100010;
        mem[9947] = 12'b000000100001;
        mem[9948] = 12'b000000100000;
        mem[9949] = 12'b000000100000;
        mem[9950] = 12'b000000011111;
        mem[9951] = 12'b000000011110;
        mem[9952] = 12'b000000011110;
        mem[9953] = 12'b000000011101;
        mem[9954] = 12'b000000011100;
        mem[9955] = 12'b000000011100;
        mem[9956] = 12'b000000011011;
        mem[9957] = 12'b000000011011;
        mem[9958] = 12'b000000011010;
        mem[9959] = 12'b000000011001;
        mem[9960] = 12'b000000011001;
        mem[9961] = 12'b000000011000;
        mem[9962] = 12'b000000010111;
        mem[9963] = 12'b000000010111;
        mem[9964] = 12'b000000010110;
        mem[9965] = 12'b000000010101;
        mem[9966] = 12'b000000010101;
        mem[9967] = 12'b000000010100;
        mem[9968] = 12'b000000010011;
        mem[9969] = 12'b000000010011;
        mem[9970] = 12'b000000010010;
        mem[9971] = 12'b000000010010;
        mem[9972] = 12'b000000010001;
        mem[9973] = 12'b000000010000;
        mem[9974] = 12'b000000010000;
        mem[9975] = 12'b000000001111;
        mem[9976] = 12'b000000001110;
        mem[9977] = 12'b000000001110;
        mem[9978] = 12'b000000001101;
        mem[9979] = 12'b000000001100;
        mem[9980] = 12'b000000001100;
        mem[9981] = 12'b000000001011;
        mem[9982] = 12'b000000001010;
        mem[9983] = 12'b000000001010;
        mem[9984] = 12'b000000001001;
        mem[9985] = 12'b000000001001;
        mem[9986] = 12'b000000001000;
        mem[9987] = 12'b000000000111;
        mem[9988] = 12'b000000000111;
        mem[9989] = 12'b000000000110;
        mem[9990] = 12'b000000000101;
        mem[9991] = 12'b000000000101;
        mem[9992] = 12'b000000000100;
        mem[9993] = 12'b000000000011;
        mem[9994] = 12'b000000000011;
        mem[9995] = 12'b000000000010;
        mem[9996] = 12'b000000000001;
        mem[9997] = 12'b000000000001;
        mem[9998] = 12'b000000000000;
        mem[9999] = 12'b000000000000;
    end

    always @(*) begin
        data1 = mem[addr1];
        data2 = mem[addr2];
        data3 = mem[addr3];
    end
endmodule
